`timescale 1ns/1ns

module sim_a_tb();


   reg 	 CLK;
   reg 	 RESET_X;
   reg 	 WR;
   reg 	 RD;
   reg [17:0] ADR;
   reg [31:0] WDATA;
   wire [31:0] RDATA;
   

   


   // clkの生成
   parameter PERIOD = 10.0; 
   
   always # (PERIOD/2) CLK = ~CLK;
   softmax_top U0 
     (
      .CLK(CLK),
      .RESET_X(RESET_X),
      .WR(WR),
      .RD(RD),
      .ADR(ADR),
      .WDATA(WDATA),
      .RDATA(RDATA)   
   );


   initial begin
      #1 CLK = 0;
     
   end

   integer i;
   integer adr_top;
   

   initial begin
      #1 RESET_X = 1; ADR = 0; WR = 0; RD = 0; WDATA = 0;
      #(PERIOD * 2) RESET_X = 0;
      #(PERIOD * 5) RESET_X = 1;

      //W0
      write(32'h00000000, 0);
      write(32'h00000004, 0);
      write(32'h00000008, 0);
      write(32'h0000000C, 0);
      write(32'h00000010, 0);
      write(32'h00000014, 0);
      write(32'h00000018, 0);
      write(32'h0000001C, 0);
      write(32'h00000020, 1);
      write(32'h00000024, 1);
      write(32'h00000028, 0);
      write(32'h0000002C, 0);
      write(32'h00000030, 0);
      write(32'h00000034, 0);
      write(32'h00000038, 0);
      write(32'h0000003C, 0);
      write(32'h00000040, 0);
      write(32'h00000044, 0);
      write(32'h00000048, 0);
      write(32'h0000004C, 0);
      write(32'h00000050, 0);
      write(32'h00000054, 0);
      write(32'h00000058, 0);
      write(32'h0000005C, 0);
      write(32'h00000060, 0);
      write(32'h00000064, 0);
      write(32'h00000068, 0);
      write(32'h0000006C, 0);
      write(32'h00000070, 0);
      write(32'h00000074, 0);
      write(32'h00000078, 0);
      write(32'h0000007C, 0);
      write(32'h00000080, 0);
      write(32'h00000084, 0);
      write(32'h00000088, -1);
      write(32'h0000008C, -1);
      write(32'h00000090, 5);
      write(32'h00000094, 10);
      write(32'h00000098, 0);
      write(32'h0000009C, -2);
      write(32'h000000A0, -2);
      write(32'h000000A4, -3);
      write(32'h000000A8, -1);
      write(32'h000000AC, 0);
      write(32'h000000B0, -1);
      write(32'h000000B4, 0);
      write(32'h000000B8, 0);
      write(32'h000000BC, -1);
      write(32'h000000C0, 0);
      write(32'h000000C4, 0);
      write(32'h000000C8, 0);
      write(32'h000000CC, 0);
      write(32'h000000D0, 0);
      write(32'h000000D4, 0);
      write(32'h000000D8, 0);
      write(32'h000000DC, 0);
      write(32'h000000E0, 0);
      write(32'h000000E4, 0);
      write(32'h000000E8, 0);
      write(32'h000000EC, -1);
      write(32'h000000F0, -2);
      write(32'h000000F4, 0);
      write(32'h000000F8, 3);
      write(32'h000000FC, -2);
      write(32'h00000100, 1);
      write(32'h00000104, 11);
      write(32'h00000108, 5);
      write(32'h0000010C, -1);
      write(32'h00000110, -8);
      write(32'h00000114, -9);
      write(32'h00000118, -3);
      write(32'h0000011C, -1);
      write(32'h00000120, 0);
      write(32'h00000124, 0);
      write(32'h00000128, 0);
      write(32'h0000012C, 0);
      write(32'h00000130, -1);
      write(32'h00000134, 0);
      write(32'h00000138, 0);
      write(32'h0000013C, 0);
      write(32'h00000140, 0);
      write(32'h00000144, 0);
      write(32'h00000148, 0);
      write(32'h0000014C, 0);
      write(32'h00000150, 0);
      write(32'h00000154, 0);
      write(32'h00000158, 1);
      write(32'h0000015C, 0);
      write(32'h00000160, -1);
      write(32'h00000164, 2);
      write(32'h00000168, 6);
      write(32'h0000016C, -1);
      write(32'h00000170, -2);
      write(32'h00000174, 5);
      write(32'h00000178, 8);
      write(32'h0000017C, 11);
      write(32'h00000180, 8);
      write(32'h00000184, -2);
      write(32'h00000188, 0);
      write(32'h0000018C, 0);
      write(32'h00000190, 1);
      write(32'h00000194, 0);
      write(32'h00000198, 2);
      write(32'h0000019C, 5);
      write(32'h000001A0, 1);
      write(32'h000001A4, -1);
      write(32'h000001A8, 0);
      write(32'h000001AC, 0);
      write(32'h000001B0, 0);
      write(32'h000001B4, 0);
      write(32'h000001B8, 0);
      write(32'h000001BC, 0);
      write(32'h000001C0, 0);
      write(32'h000001C4, 1);
      write(32'h000001C8, 4);
      write(32'h000001CC, 0);
      write(32'h000001D0, -2);
      write(32'h000001D4, -1);
      write(32'h000001D8, 5);
      write(32'h000001DC, 0);
      write(32'h000001E0, -5);
      write(32'h000001E4, 2);
      write(32'h000001E8, 6);
      write(32'h000001EC, 7);
      write(32'h000001F0, 0);
      write(32'h000001F4, 0);
      write(32'h000001F8, 8);
      write(32'h000001FC, -3);
      write(32'h00000200, -3);
      write(32'h00000204, -5);
      write(32'h00000208, -1);
      write(32'h0000020C, 6);
      write(32'h00000210, 0);
      write(32'h00000214, -2);
      write(32'h00000218, 0);
      write(32'h0000021C, 0);
      write(32'h00000220, 0);
      write(32'h00000224, 0);
      write(32'h00000228, 0);
      write(32'h0000022C, 0);
      write(32'h00000230, 0);
      write(32'h00000234, 2);
      write(32'h00000238, 0);
      write(32'h0000023C, -1);
      write(32'h00000240, 0);
      write(32'h00000244, 0);
      write(32'h00000248, 0);
      write(32'h0000024C, 5);
      write(32'h00000250, 10);
      write(32'h00000254, 20);
      write(32'h00000258, 13);
      write(32'h0000025C, 4);
      write(32'h00000260, 0);
      write(32'h00000264, 4);
      write(32'h00000268, 20);
      write(32'h0000026C, 5);
      write(32'h00000270, -5);
      write(32'h00000274, -8);
      write(32'h00000278, -8);
      write(32'h0000027C, -3);
      write(32'h00000280, 0);
      write(32'h00000284, 0);
      write(32'h00000288, -1);
      write(32'h0000028C, 0);
      write(32'h00000290, 0);
      write(32'h00000294, 0);
      write(32'h00000298, 0);
      write(32'h0000029C, 0);
      write(32'h000002A0, 0);
      write(32'h000002A4, 0);
      write(32'h000002A8, -1);
      write(32'h000002AC, 6);
      write(32'h000002B0, 4);
      write(32'h000002B4, 5);
      write(32'h000002B8, 1);
      write(32'h000002BC, 2);
      write(32'h000002C0, 21);
      write(32'h000002C4, 28);
      write(32'h000002C8, 11);
      write(32'h000002CC, -2);
      write(32'h000002D0, -14);
      write(32'h000002D4, -13);
      write(32'h000002D8, -4);
      write(32'h000002DC, -9);
      write(32'h000002E0, -20);
      write(32'h000002E4, -18);
      write(32'h000002E8, -12);
      write(32'h000002EC, -14);
      write(32'h000002F0, -8);
      write(32'h000002F4, -1);
      write(32'h000002F8, -1);
      write(32'h000002FC, 0);
      write(32'h00000300, 0);
      write(32'h00000304, 0);
      write(32'h00000308, 0);
      write(32'h0000030C, 0);
      write(32'h00000310, 0);
      write(32'h00000314, 0);
      write(32'h00000318, 0);
      write(32'h0000031C, 7);
      write(32'h00000320, 4);
      write(32'h00000324, 0);
      write(32'h00000328, 0);
      write(32'h0000032C, 5);
      write(32'h00000330, 10);
      write(32'h00000334, 17);
      write(32'h00000338, -1);
      write(32'h0000033C, -15);
      write(32'h00000340, -16);
      write(32'h00000344, -8);
      write(32'h00000348, -3);
      write(32'h0000034C, -2);
      write(32'h00000350, -3);
      write(32'h00000354, -4);
      write(32'h00000358, -2);
      write(32'h0000035C, -6);
      write(32'h00000360, -3);
      write(32'h00000364, -3);
      write(32'h00000368, -4);
      write(32'h0000036C, 0);
      write(32'h00000370, 0);
      write(32'h00000374, 0);
      write(32'h00000378, 0);
      write(32'h0000037C, 0);
      write(32'h00000380, 0);
      write(32'h00000384, 0);
      write(32'h00000388, -2);
      write(32'h0000038C, 0);
      write(32'h00000390, 0);
      write(32'h00000394, -3);
      write(32'h00000398, 2);
      write(32'h0000039C, 0);
      write(32'h000003A0, -1);
      write(32'h000003A4, 7);
      write(32'h000003A8, 2);
      write(32'h000003AC, -5);
      write(32'h000003B0, -4);
      write(32'h000003B4, 7);
      write(32'h000003B8, 3);
      write(32'h000003BC, 1);
      write(32'h000003C0, 5);
      write(32'h000003C4, 5);
      write(32'h000003C8, -5);
      write(32'h000003CC, -6);
      write(32'h000003D0, -4);
      write(32'h000003D4, -5);
      write(32'h000003D8, -6);
      write(32'h000003DC, 0);
      write(32'h000003E0, 0);
      write(32'h000003E4, 0);
      write(32'h000003E8, 0);
      write(32'h000003EC, 0);
      write(32'h000003F0, 0);
      write(32'h000003F4, 0);
      write(32'h000003F8, 1);
      write(32'h000003FC, -5);
      write(32'h00000400, -8);
      write(32'h00000404, -16);
      write(32'h00000408, -2);
      write(32'h0000040C, 2);
      write(32'h00000410, -2);
      write(32'h00000414, 12);
      write(32'h00000418, 5);
      write(32'h0000041C, -1);
      write(32'h00000420, -2);
      write(32'h00000424, 1);
      write(32'h00000428, 6);
      write(32'h0000042C, 9);
      write(32'h00000430, 13);
      write(32'h00000434, 9);
      write(32'h00000438, -6);
      write(32'h0000043C, -13);
      write(32'h00000440, -14);
      write(32'h00000444, -12);
      write(32'h00000448, -4);
      write(32'h0000044C, 0);
      write(32'h00000450, 0);
      write(32'h00000454, 0);
      write(32'h00000458, 0);
      write(32'h0000045C, 0);
      write(32'h00000460, 0);
      write(32'h00000464, 0);
      write(32'h00000468, -4);
      write(32'h0000046C, -14);
      write(32'h00000470, -15);
      write(32'h00000474, -15);
      write(32'h00000478, -6);
      write(32'h0000047C, -7);
      write(32'h00000480, -1);
      write(32'h00000484, 10);
      write(32'h00000488, 5);
      write(32'h0000048C, 8);
      write(32'h00000490, 1);
      write(32'h00000494, 5);
      write(32'h00000498, 15);
      write(32'h0000049C, 12);
      write(32'h000004A0, 8);
      write(32'h000004A4, 17);
      write(32'h000004A8, 3);
      write(32'h000004AC, -5);
      write(32'h000004B0, -10);
      write(32'h000004B4, -11);
      write(32'h000004B8, -6);
      write(32'h000004BC, 0);
      write(32'h000004C0, 0);
      write(32'h000004C4, 0);
      write(32'h000004C8, 0);
      write(32'h000004CC, 0);
      write(32'h000004D0, 0);
      write(32'h000004D4, -1);
      write(32'h000004D8, -6);
      write(32'h000004DC, -16);
      write(32'h000004E0, -9);
      write(32'h000004E4, -1);
      write(32'h000004E8, -9);
      write(32'h000004EC, -15);
      write(32'h000004F0, 9);
      write(32'h000004F4, 10);
      write(32'h000004F8, -3);
      write(32'h000004FC, -1);
      write(32'h00000500, -2);
      write(32'h00000504, 1);
      write(32'h00000508, 3);
      write(32'h0000050C, 3);
      write(32'h00000510, 2);
      write(32'h00000514, 5);
      write(32'h00000518, 6);
      write(32'h0000051C, -7);
      write(32'h00000520, -8);
      write(32'h00000524, -7);
      write(32'h00000528, -8);
      write(32'h0000052C, -2);
      write(32'h00000530, 0);
      write(32'h00000534, 0);
      write(32'h00000538, 0);
      write(32'h0000053C, 0);
      write(32'h00000540, 0);
      write(32'h00000544, 0);
      write(32'h00000548, -3);
      write(32'h0000054C, -3);
      write(32'h00000550, -1);
      write(32'h00000554, -12);
      write(32'h00000558, -20);
      write(32'h0000055C, -5);
      write(32'h00000560, 18);
      write(32'h00000564, 5);
      write(32'h00000568, -1);
      write(32'h0000056C, -7);
      write(32'h00000570, -4);
      write(32'h00000574, 11);
      write(32'h00000578, 7);
      write(32'h0000057C, 2);
      write(32'h00000580, 6);
      write(32'h00000584, 7);
      write(32'h00000588, 8);
      write(32'h0000058C, 0);
      write(32'h00000590, -7);
      write(32'h00000594, -2);
      write(32'h00000598, -3);
      write(32'h0000059C, -1);
      write(32'h000005A0, 0);
      write(32'h000005A4, 0);
      write(32'h000005A8, 0);
      write(32'h000005AC, 0);
      write(32'h000005B0, 0);
      write(32'h000005B4, 0);
      write(32'h000005B8, 0);
      write(32'h000005BC, 0);
      write(32'h000005C0, -9);
      write(32'h000005C4, -19);
      write(32'h000005C8, -11);
      write(32'h000005CC, 3);
      write(32'h000005D0, 10);
      write(32'h000005D4, 6);
      write(32'h000005D8, -5);
      write(32'h000005DC, -18);
      write(32'h000005E0, -6);
      write(32'h000005E4, 9);
      write(32'h000005E8, 14);
      write(32'h000005EC, 15);
      write(32'h000005F0, 5);
      write(32'h000005F4, -8);
      write(32'h000005F8, 6);
      write(32'h000005FC, 10);
      write(32'h00000600, -4);
      write(32'h00000604, -2);
      write(32'h00000608, 1);
      write(32'h0000060C, 0);
      write(32'h00000610, 0);
      write(32'h00000614, 0);
      write(32'h00000618, 0);
      write(32'h0000061C, 0);
      write(32'h00000620, 0);
      write(32'h00000624, 1);
      write(32'h00000628, 0);
      write(32'h0000062C, -1);
      write(32'h00000630, -9);
      write(32'h00000634, -2);
      write(32'h00000638, 1);
      write(32'h0000063C, 2);
      write(32'h00000640, 4);
      write(32'h00000644, 25);
      write(32'h00000648, 6);
      write(32'h0000064C, 6);
      write(32'h00000650, 11);
      write(32'h00000654, 3);
      write(32'h00000658, 8);
      write(32'h0000065C, 14);
      write(32'h00000660, -6);
      write(32'h00000664, -12);
      write(32'h00000668, 3);
      write(32'h0000066C, 15);
      write(32'h00000670, 5);
      write(32'h00000674, 0);
      write(32'h00000678, 5);
      write(32'h0000067C, 0);
      write(32'h00000680, 0);
      write(32'h00000684, 0);
      write(32'h00000688, 0);
      write(32'h0000068C, 0);
      write(32'h00000690, 0);
      write(32'h00000694, 3);
      write(32'h00000698, 1);
      write(32'h0000069C, 0);
      write(32'h000006A0, 3);
      write(32'h000006A4, 9);
      write(32'h000006A8, 3);
      write(32'h000006AC, -11);
      write(32'h000006B0, 1);
      write(32'h000006B4, 25);
      write(32'h000006B8, 21);
      write(32'h000006BC, 19);
      write(32'h000006C0, 5);
      write(32'h000006C4, -3);
      write(32'h000006C8, -2);
      write(32'h000006CC, -1);
      write(32'h000006D0, -12);
      write(32'h000006D4, -5);
      write(32'h000006D8, 5);
      write(32'h000006DC, 12);
      write(32'h000006E0, 12);
      write(32'h000006E4, 8);
      write(32'h000006E8, 4);
      write(32'h000006EC, 0);
      write(32'h000006F0, 0);
      write(32'h000006F4, 0);
      write(32'h000006F8, 0);
      write(32'h000006FC, 0);
      write(32'h00000700, 0);
      write(32'h00000704, 4);
      write(32'h00000708, 0);
      write(32'h0000070C, 7);
      write(32'h00000710, 8);
      write(32'h00000714, 8);
      write(32'h00000718, 0);
      write(32'h0000071C, -14);
      write(32'h00000720, -4);
      write(32'h00000724, 21);
      write(32'h00000728, 30);
      write(32'h0000072C, 10);
      write(32'h00000730, -3);
      write(32'h00000734, -7);
      write(32'h00000738, 0);
      write(32'h0000073C, -11);
      write(32'h00000740, -21);
      write(32'h00000744, -7);
      write(32'h00000748, 10);
      write(32'h0000074C, 11);
      write(32'h00000750, 9);
      write(32'h00000754, 10);
      write(32'h00000758, 4);
      write(32'h0000075C, 0);
      write(32'h00000760, 0);
      write(32'h00000764, 0);
      write(32'h00000768, 0);
      write(32'h0000076C, 0);
      write(32'h00000770, 0);
      write(32'h00000774, 5);
      write(32'h00000778, 2);
      write(32'h0000077C, 9);
      write(32'h00000780, 3);
      write(32'h00000784, 7);
      write(32'h00000788, 2);
      write(32'h0000078C, -14);
      write(32'h00000790, 2);
      write(32'h00000794, 15);
      write(32'h00000798, 29);
      write(32'h0000079C, 6);
      write(32'h000007A0, -9);
      write(32'h000007A4, 6);
      write(32'h000007A8, 12);
      write(32'h000007AC, -16);
      write(32'h000007B0, -21);
      write(32'h000007B4, -4);
      write(32'h000007B8, 1);
      write(32'h000007BC, 6);
      write(32'h000007C0, 15);
      write(32'h000007C4, 10);
      write(32'h000007C8, 3);
      write(32'h000007CC, 0);
      write(32'h000007D0, 0);
      write(32'h000007D4, 0);
      write(32'h000007D8, 0);
      write(32'h000007DC, 0);
      write(32'h000007E0, 0);
      write(32'h000007E4, 3);
      write(32'h000007E8, 7);
      write(32'h000007EC, 6);
      write(32'h000007F0, 5);
      write(32'h000007F4, 14);
      write(32'h000007F8, 14);
      write(32'h000007FC, 5);
      write(32'h00000800, 0);
      write(32'h00000804, 0);
      write(32'h00000808, 24);
      write(32'h0000080C, 13);
      write(32'h00000810, -2);
      write(32'h00000814, 1);
      write(32'h00000818, -5);
      write(32'h0000081C, -8);
      write(32'h00000820, -3);
      write(32'h00000824, -5);
      write(32'h00000828, -7);
      write(32'h0000082C, -2);
      write(32'h00000830, 11);
      write(32'h00000834, 10);
      write(32'h00000838, 4);
      write(32'h0000083C, 0);
      write(32'h00000840, 0);
      write(32'h00000844, 0);
      write(32'h00000848, 0);
      write(32'h0000084C, 0);
      write(32'h00000850, 0);
      write(32'h00000854, 1);
      write(32'h00000858, 7);
      write(32'h0000085C, 12);
      write(32'h00000860, 9);
      write(32'h00000864, 7);
      write(32'h00000868, 13);
      write(32'h0000086C, -2);
      write(32'h00000870, -15);
      write(32'h00000874, -8);
      write(32'h00000878, 4);
      write(32'h0000087C, 4);
      write(32'h00000880, 3);
      write(32'h00000884, -4);
      write(32'h00000888, -15);
      write(32'h0000088C, -2);
      write(32'h00000890, 10);
      write(32'h00000894, 4);
      write(32'h00000898, -2);
      write(32'h0000089C, -2);
      write(32'h000008A0, 0);
      write(32'h000008A4, 7);
      write(32'h000008A8, 3);
      write(32'h000008AC, 0);
      write(32'h000008B0, 0);
      write(32'h000008B4, 0);
      write(32'h000008B8, 0);
      write(32'h000008BC, 0);
      write(32'h000008C0, 0);
      write(32'h000008C4, 2);
      write(32'h000008C8, 3);
      write(32'h000008CC, 10);
      write(32'h000008D0, 11);
      write(32'h000008D4, 3);
      write(32'h000008D8, 1);
      write(32'h000008DC, -3);
      write(32'h000008E0, -5);
      write(32'h000008E4, 5);
      write(32'h000008E8, 1);
      write(32'h000008EC, 2);
      write(32'h000008F0, -8);
      write(32'h000008F4, -8);
      write(32'h000008F8, -1);
      write(32'h000008FC, -3);
      write(32'h00000900, -2);
      write(32'h00000904, 0);
      write(32'h00000908, 7);
      write(32'h0000090C, -7);
      write(32'h00000910, -4);
      write(32'h00000914, 5);
      write(32'h00000918, 3);
      write(32'h0000091C, 0);
      write(32'h00000920, 0);
      write(32'h00000924, 0);
      write(32'h00000928, 0);
      write(32'h0000092C, 0);
      write(32'h00000930, 0);
      write(32'h00000934, 2);
      write(32'h00000938, 3);
      write(32'h0000093C, 6);
      write(32'h00000940, -3);
      write(32'h00000944, -6);
      write(32'h00000948, 0);
      write(32'h0000094C, 0);
      write(32'h00000950, -5);
      write(32'h00000954, 0);
      write(32'h00000958, 5);
      write(32'h0000095C, 9);
      write(32'h00000960, -5);
      write(32'h00000964, 14);
      write(32'h00000968, 5);
      write(32'h0000096C, -8);
      write(32'h00000970, -5);
      write(32'h00000974, -10);
      write(32'h00000978, -6);
      write(32'h0000097C, -2);
      write(32'h00000980, 2);
      write(32'h00000984, 4);
      write(32'h00000988, 3);
      write(32'h0000098C, 0);
      write(32'h00000990, 0);
      write(32'h00000994, 0);
      write(32'h00000998, 0);
      write(32'h0000099C, 0);
      write(32'h000009A0, 0);
      write(32'h000009A4, 2);
      write(32'h000009A8, 2);
      write(32'h000009AC, 8);
      write(32'h000009B0, -2);
      write(32'h000009B4, -4);
      write(32'h000009B8, 4);
      write(32'h000009BC, 2);
      write(32'h000009C0, -11);
      write(32'h000009C4, -4);
      write(32'h000009C8, 12);
      write(32'h000009CC, 11);
      write(32'h000009D0, 3);
      write(32'h000009D4, 11);
      write(32'h000009D8, -3);
      write(32'h000009DC, -9);
      write(32'h000009E0, -12);
      write(32'h000009E4, -5);
      write(32'h000009E8, -1);
      write(32'h000009EC, 8);
      write(32'h000009F0, 4);
      write(32'h000009F4, 4);
      write(32'h000009F8, 1);
      write(32'h000009FC, 0);
      write(32'h00000A00, 0);
      write(32'h00000A04, 0);
      write(32'h00000A08, 0);
      write(32'h00000A0C, 0);
      write(32'h00000A10, 0);
      write(32'h00000A14, 1);
      write(32'h00000A18, 2);
      write(32'h00000A1C, 7);
      write(32'h00000A20, 3);
      write(32'h00000A24, 6);
      write(32'h00000A28, 8);
      write(32'h00000A2C, -1);
      write(32'h00000A30, -8);
      write(32'h00000A34, -2);
      write(32'h00000A38, 4);
      write(32'h00000A3C, 10);
      write(32'h00000A40, 7);
      write(32'h00000A44, -6);
      write(32'h00000A48, -17);
      write(32'h00000A4C, -12);
      write(32'h00000A50, -9);
      write(32'h00000A54, 0);
      write(32'h00000A58, 3);
      write(32'h00000A5C, 13);
      write(32'h00000A60, 2);
      write(32'h00000A64, 0);
      write(32'h00000A68, -1);
      write(32'h00000A6C, 0);
      write(32'h00000A70, 0);
      write(32'h00000A74, 0);
      write(32'h00000A78, 0);
      write(32'h00000A7C, 0);
      write(32'h00000A80, 0);
      write(32'h00000A84, 0);
      write(32'h00000A88, 1);
      write(32'h00000A8C, 7);
      write(32'h00000A90, 13);
      write(32'h00000A94, 12);
      write(32'h00000A98, 5);
      write(32'h00000A9C, -6);
      write(32'h00000AA0, -5);
      write(32'h00000AA4, -9);
      write(32'h00000AA8, -1);
      write(32'h00000AAC, 11);
      write(32'h00000AB0, 0);
      write(32'h00000AB4, -19);
      write(32'h00000AB8, -20);
      write(32'h00000ABC, -8);
      write(32'h00000AC0, -2);
      write(32'h00000AC4, 6);
      write(32'h00000AC8, 7);
      write(32'h00000ACC, 8);
      write(32'h00000AD0, -2);
      write(32'h00000AD4, -3);
      write(32'h00000AD8, -1);
      write(32'h00000ADC, 0);
      write(32'h00000AE0, 0);
      write(32'h00000AE4, 0);
      write(32'h00000AE8, 0);
      write(32'h00000AEC, 0);
      write(32'h00000AF0, 0);
      write(32'h00000AF4, 0);
      write(32'h00000AF8, -1);
      write(32'h00000AFC, 1);
      write(32'h00000B00, 12);
      write(32'h00000B04, 18);
      write(32'h00000B08, 8);
      write(32'h00000B0C, -2);
      write(32'h00000B10, -6);
      write(32'h00000B14, -11);
      write(32'h00000B18, -2);
      write(32'h00000B1C, 4);
      write(32'h00000B20, -6);
      write(32'h00000B24, -18);
      write(32'h00000B28, -11);
      write(32'h00000B2C, -5);
      write(32'h00000B30, 1);
      write(32'h00000B34, 0);
      write(32'h00000B38, 1);
      write(32'h00000B3C, 1);
      write(32'h00000B40, -4);
      write(32'h00000B44, -2);
      write(32'h00000B48, 0);
      write(32'h00000B4C, 0);
      write(32'h00000B50, 0);
      write(32'h00000B54, 0);
      write(32'h00000B58, 0);
      write(32'h00000B5C, 0);
      write(32'h00000B60, 0);
      write(32'h00000B64, 0);
      write(32'h00000B68, 0);
      write(32'h00000B6C, -1);
      write(32'h00000B70, 7);
      write(32'h00000B74, 11);
      write(32'h00000B78, 7);
      write(32'h00000B7C, 4);
      write(32'h00000B80, 3);
      write(32'h00000B84, 0);
      write(32'h00000B88, 2);
      write(32'h00000B8C, 7);
      write(32'h00000B90, -1);
      write(32'h00000B94, -14);
      write(32'h00000B98, -4);
      write(32'h00000B9C, 0);
      write(32'h00000BA0, -4);
      write(32'h00000BA4, -2);
      write(32'h00000BA8, 3);
      write(32'h00000BAC, 0);
      write(32'h00000BB0, -2);
      write(32'h00000BB4, 0);
      write(32'h00000BB8, 0);
      write(32'h00000BBC, 0);
      write(32'h00000BC0, 0);
      write(32'h00000BC4, 0);
      write(32'h00000BC8, 0);
      write(32'h00000BCC, 0);
      write(32'h00000BD0, 0);
      write(32'h00000BD4, 0);
      write(32'h00000BD8, 0);
      write(32'h00000BDC, 0);
      write(32'h00000BE0, 4);
      write(32'h00000BE4, 14);
      write(32'h00000BE8, 12);
      write(32'h00000BEC, 8);
      write(32'h00000BF0, 3);
      write(32'h00000BF4, -7);
      write(32'h00000BF8, -6);
      write(32'h00000BFC, -2);
      write(32'h00000C00, -10);
      write(32'h00000C04, -9);
      write(32'h00000C08, -4);
      write(32'h00000C0C, -3);
      write(32'h00000C10, 1);
      write(32'h00000C14, 5);
      write(32'h00000C18, 1);
      write(32'h00000C1C, -1);
      write(32'h00000C20, 0);
      write(32'h00000C24, 0);
      write(32'h00000C28, 0);
      write(32'h00000C2C, 0);
      write(32'h00000C30, 0);
      write(32'h00000C34, 0);
      write(32'h00000C38, 0);
      write(32'h00000C3C, 0);

      #(PERIOD * 20) ;
      
      //W1
      write(32'h00001000, 0);
      write(32'h00001004, 0);
      write(32'h00001008, 0);
      write(32'h0000100C, 0);
      write(32'h00001010, 0);
      write(32'h00001014, 0);
      write(32'h00001018, 0);
      write(32'h0000101C, 0);
      write(32'h00001020, 0);
      write(32'h00001024, 0);
      write(32'h00001028, 0);
      write(32'h0000102C, 0);
      write(32'h00001030, 0);
      write(32'h00001034, 0);
      write(32'h00001038, 0);
      write(32'h0000103C, 0);
      write(32'h00001040, 0);
      write(32'h00001044, 0);
      write(32'h00001048, 0);
      write(32'h0000104C, 0);
      write(32'h00001050, 0);
      write(32'h00001054, 0);
      write(32'h00001058, 0);
      write(32'h0000105C, 0);
      write(32'h00001060, 0);
      write(32'h00001064, 0);
      write(32'h00001068, 0);
      write(32'h0000106C, 0);
      write(32'h00001070, 0);
      write(32'h00001074, 0);
      write(32'h00001078, 0);
      write(32'h0000107C, 0);
      write(32'h00001080, 0);
      write(32'h00001084, 0);
      write(32'h00001088, -1);
      write(32'h0000108C, 0);
      write(32'h00001090, 0);
      write(32'h00001094, 0);
      write(32'h00001098, 0);
      write(32'h0000109C, 0);
      write(32'h000010A0, 0);
      write(32'h000010A4, 0);
      write(32'h000010A8, 0);
      write(32'h000010AC, 0);
      write(32'h000010B0, 0);
      write(32'h000010B4, 0);
      write(32'h000010B8, 0);
      write(32'h000010BC, 0);
      write(32'h000010C0, 0);
      write(32'h000010C4, 0);
      write(32'h000010C8, 0);
      write(32'h000010CC, 0);
      write(32'h000010D0, 0);
      write(32'h000010D4, 0);
      write(32'h000010D8, 0);
      write(32'h000010DC, 0);
      write(32'h000010E0, 0);
      write(32'h000010E4, 0);
      write(32'h000010E8, 0);
      write(32'h000010EC, 0);
      write(32'h000010F0, -2);
      write(32'h000010F4, -2);
      write(32'h000010F8, -2);
      write(32'h000010FC, -1);
      write(32'h00001100, -1);
      write(32'h00001104, -2);
      write(32'h00001108, -2);
      write(32'h0000110C, -1);
      write(32'h00001110, -1);
      write(32'h00001114, -1);
      write(32'h00001118, -1);
      write(32'h0000111C, -1);
      write(32'h00001120, -1);
      write(32'h00001124, 0);
      write(32'h00001128, 0);
      write(32'h0000112C, 0);
      write(32'h00001130, 0);
      write(32'h00001134, 0);
      write(32'h00001138, 0);
      write(32'h0000113C, 0);
      write(32'h00001140, 0);
      write(32'h00001144, 0);
      write(32'h00001148, 0);
      write(32'h0000114C, 0);
      write(32'h00001150, 0);
      write(32'h00001154, 0);
      write(32'h00001158, 1);
      write(32'h0000115C, 1);
      write(32'h00001160, -1);
      write(32'h00001164, -2);
      write(32'h00001168, -5);
      write(32'h0000116C, -5);
      write(32'h00001170, -3);
      write(32'h00001174, -3);
      write(32'h00001178, -3);
      write(32'h0000117C, -3);
      write(32'h00001180, -3);
      write(32'h00001184, -3);
      write(32'h00001188, -3);
      write(32'h0000118C, -3);
      write(32'h00001190, -5);
      write(32'h00001194, -7);
      write(32'h00001198, -3);
      write(32'h0000119C, 0);
      write(32'h000011A0, 0);
      write(32'h000011A4, 0);
      write(32'h000011A8, 0);
      write(32'h000011AC, 0);
      write(32'h000011B0, 0);
      write(32'h000011B4, 0);
      write(32'h000011B8, 0);
      write(32'h000011BC, 0);
      write(32'h000011C0, 0);
      write(32'h000011C4, 1);
      write(32'h000011C8, 9);
      write(32'h000011CC, 7);
      write(32'h000011D0, 1);
      write(32'h000011D4, -1);
      write(32'h000011D8, -8);
      write(32'h000011DC, -10);
      write(32'h000011E0, -9);
      write(32'h000011E4, -5);
      write(32'h000011E8, -5);
      write(32'h000011EC, -4);
      write(32'h000011F0, -4);
      write(32'h000011F4, -4);
      write(32'h000011F8, -4);
      write(32'h000011FC, -5);
      write(32'h00001200, -8);
      write(32'h00001204, -9);
      write(32'h00001208, -9);
      write(32'h0000120C, -2);
      write(32'h00001210, 0);
      write(32'h00001214, 0);
      write(32'h00001218, 0);
      write(32'h0000121C, 0);
      write(32'h00001220, 0);
      write(32'h00001224, 0);
      write(32'h00001228, 0);
      write(32'h0000122C, 0);
      write(32'h00001230, 0);
      write(32'h00001234, 1);
      write(32'h00001238, 7);
      write(32'h0000123C, 15);
      write(32'h00001240, 8);
      write(32'h00001244, -4);
      write(32'h00001248, -4);
      write(32'h0000124C, -11);
      write(32'h00001250, -9);
      write(32'h00001254, -6);
      write(32'h00001258, -6);
      write(32'h0000125C, -7);
      write(32'h00001260, -7);
      write(32'h00001264, -6);
      write(32'h00001268, -5);
      write(32'h0000126C, -4);
      write(32'h00001270, -3);
      write(32'h00001274, -4);
      write(32'h00001278, -7);
      write(32'h0000127C, -5);
      write(32'h00001280, 0);
      write(32'h00001284, 0);
      write(32'h00001288, 0);
      write(32'h0000128C, 0);
      write(32'h00001290, 0);
      write(32'h00001294, 0);
      write(32'h00001298, 0);
      write(32'h0000129C, 0);
      write(32'h000012A0, 0);
      write(32'h000012A4, 1);
      write(32'h000012A8, 5);
      write(32'h000012AC, 11);
      write(32'h000012B0, 13);
      write(32'h000012B4, -1);
      write(32'h000012B8, -6);
      write(32'h000012BC, -13);
      write(32'h000012C0, -10);
      write(32'h000012C4, -10);
      write(32'h000012C8, -10);
      write(32'h000012CC, -10);
      write(32'h000012D0, -8);
      write(32'h000012D4, -7);
      write(32'h000012D8, -6);
      write(32'h000012DC, -2);
      write(32'h000012E0, -3);
      write(32'h000012E4, 1);
      write(32'h000012E8, -3);
      write(32'h000012EC, -6);
      write(32'h000012F0, -1);
      write(32'h000012F4, 0);
      write(32'h000012F8, 0);
      write(32'h000012FC, 0);
      write(32'h00001300, 0);
      write(32'h00001304, 0);
      write(32'h00001308, 0);
      write(32'h0000130C, 0);
      write(32'h00001310, 0);
      write(32'h00001314, 1);
      write(32'h00001318, 6);
      write(32'h0000131C, 10);
      write(32'h00001320, 14);
      write(32'h00001324, 6);
      write(32'h00001328, -8);
      write(32'h0000132C, -14);
      write(32'h00001330, -12);
      write(32'h00001334, -12);
      write(32'h00001338, -10);
      write(32'h0000133C, -11);
      write(32'h00001340, -10);
      write(32'h00001344, -9);
      write(32'h00001348, -8);
      write(32'h0000134C, -3);
      write(32'h00001350, 1);
      write(32'h00001354, -1);
      write(32'h00001358, 4);
      write(32'h0000135C, -3);
      write(32'h00001360, -2);
      write(32'h00001364, 0);
      write(32'h00001368, 0);
      write(32'h0000136C, 0);
      write(32'h00001370, 0);
      write(32'h00001374, 0);
      write(32'h00001378, 0);
      write(32'h0000137C, 0);
      write(32'h00001380, 0);
      write(32'h00001384, 2);
      write(32'h00001388, 7);
      write(32'h0000138C, 10);
      write(32'h00001390, 16);
      write(32'h00001394, 9);
      write(32'h00001398, -11);
      write(32'h0000139C, -12);
      write(32'h000013A0, -11);
      write(32'h000013A4, -10);
      write(32'h000013A8, -9);
      write(32'h000013AC, -10);
      write(32'h000013B0, -9);
      write(32'h000013B4, -8);
      write(32'h000013B8, -8);
      write(32'h000013BC, -6);
      write(32'h000013C0, 1);
      write(32'h000013C4, 5);
      write(32'h000013C8, 4);
      write(32'h000013CC, 5);
      write(32'h000013D0, -1);
      write(32'h000013D4, 0);
      write(32'h000013D8, 0);
      write(32'h000013DC, 0);
      write(32'h000013E0, 0);
      write(32'h000013E4, 0);
      write(32'h000013E8, 0);
      write(32'h000013EC, 0);
      write(32'h000013F0, 0);
      write(32'h000013F4, 2);
      write(32'h000013F8, 6);
      write(32'h000013FC, 11);
      write(32'h00001400, 21);
      write(32'h00001404, 9);
      write(32'h00001408, -11);
      write(32'h0000140C, -10);
      write(32'h00001410, -11);
      write(32'h00001414, -9);
      write(32'h00001418, -9);
      write(32'h0000141C, -11);
      write(32'h00001420, -10);
      write(32'h00001424, -9);
      write(32'h00001428, -8);
      write(32'h0000142C, -3);
      write(32'h00001430, -1);
      write(32'h00001434, 4);
      write(32'h00001438, 9);
      write(32'h0000143C, 7);
      write(32'h00001440, 4);
      write(32'h00001444, 0);
      write(32'h00001448, 0);
      write(32'h0000144C, 0);
      write(32'h00001450, 0);
      write(32'h00001454, 0);
      write(32'h00001458, 0);
      write(32'h0000145C, 0);
      write(32'h00001460, 0);
      write(32'h00001464, 2);
      write(32'h00001468, 5);
      write(32'h0000146C, 10);
      write(32'h00001470, 21);
      write(32'h00001474, 7);
      write(32'h00001478, -10);
      write(32'h0000147C, -10);
      write(32'h00001480, -11);
      write(32'h00001484, -11);
      write(32'h00001488, -11);
      write(32'h0000148C, -11);
      write(32'h00001490, -11);
      write(32'h00001494, -11);
      write(32'h00001498, -10);
      write(32'h0000149C, -3);
      write(32'h000014A0, 5);
      write(32'h000014A4, 0);
      write(32'h000014A8, 11);
      write(32'h000014AC, 12);
      write(32'h000014B0, 7);
      write(32'h000014B4, 4);
      write(32'h000014B8, 0);
      write(32'h000014BC, 0);
      write(32'h000014C0, 0);
      write(32'h000014C4, 0);
      write(32'h000014C8, 0);
      write(32'h000014CC, 0);
      write(32'h000014D0, 0);
      write(32'h000014D4, 2);
      write(32'h000014D8, 6);
      write(32'h000014DC, 10);
      write(32'h000014E0, 21);
      write(32'h000014E4, 8);
      write(32'h000014E8, -9);
      write(32'h000014EC, -11);
      write(32'h000014F0, -11);
      write(32'h000014F4, -8);
      write(32'h000014F8, -8);
      write(32'h000014FC, -11);
      write(32'h00001500, -11);
      write(32'h00001504, -10);
      write(32'h00001508, -10);
      write(32'h0000150C, -8);
      write(32'h00001510, 2);
      write(32'h00001514, 5);
      write(32'h00001518, 7);
      write(32'h0000151C, 16);
      write(32'h00001520, 11);
      write(32'h00001524, 9);
      write(32'h00001528, 0);
      write(32'h0000152C, 0);
      write(32'h00001530, 0);
      write(32'h00001534, 0);
      write(32'h00001538, 0);
      write(32'h0000153C, 0);
      write(32'h00001540, 0);
      write(32'h00001544, 2);
      write(32'h00001548, 5);
      write(32'h0000154C, 9);
      write(32'h00001550, 18);
      write(32'h00001554, 15);
      write(32'h00001558, 2);
      write(32'h0000155C, -10);
      write(32'h00001560, -11);
      write(32'h00001564, -6);
      write(32'h00001568, -6);
      write(32'h0000156C, -9);
      write(32'h00001570, -10);
      write(32'h00001574, -9);
      write(32'h00001578, -8);
      write(32'h0000157C, -7);
      write(32'h00001580, -1);
      write(32'h00001584, 6);
      write(32'h00001588, 7);
      write(32'h0000158C, 17);
      write(32'h00001590, 17);
      write(32'h00001594, 11);
      write(32'h00001598, 1);
      write(32'h0000159C, 0);
      write(32'h000015A0, 0);
      write(32'h000015A4, 0);
      write(32'h000015A8, 0);
      write(32'h000015AC, 0);
      write(32'h000015B0, 0);
      write(32'h000015B4, 2);
      write(32'h000015B8, 4);
      write(32'h000015BC, 8);
      write(32'h000015C0, 15);
      write(32'h000015C4, 17);
      write(32'h000015C8, 11);
      write(32'h000015CC, -8);
      write(32'h000015D0, -7);
      write(32'h000015D4, -1);
      write(32'h000015D8, -1);
      write(32'h000015DC, -7);
      write(32'h000015E0, -8);
      write(32'h000015E4, -7);
      write(32'h000015E8, -6);
      write(32'h000015EC, -4);
      write(32'h000015F0, 0);
      write(32'h000015F4, 3);
      write(32'h000015F8, 9);
      write(32'h000015FC, 16);
      write(32'h00001600, 18);
      write(32'h00001604, 16);
      write(32'h00001608, 3);
      write(32'h0000160C, 0);
      write(32'h00001610, 0);
      write(32'h00001614, 0);
      write(32'h00001618, 0);
      write(32'h0000161C, 0);
      write(32'h00001620, 0);
      write(32'h00001624, 3);
      write(32'h00001628, 5);
      write(32'h0000162C, 6);
      write(32'h00001630, 14);
      write(32'h00001634, 17);
      write(32'h00001638, 13);
      write(32'h0000163C, -3);
      write(32'h00001640, 0);
      write(32'h00001644, 5);
      write(32'h00001648, 3);
      write(32'h0000164C, -6);
      write(32'h00001650, -8);
      write(32'h00001654, -8);
      write(32'h00001658, -7);
      write(32'h0000165C, 0);
      write(32'h00001660, 5);
      write(32'h00001664, 6);
      write(32'h00001668, 12);
      write(32'h0000166C, 18);
      write(32'h00001670, 14);
      write(32'h00001674, 19);
      write(32'h00001678, 2);
      write(32'h0000167C, 0);
      write(32'h00001680, 0);
      write(32'h00001684, 0);
      write(32'h00001688, 0);
      write(32'h0000168C, 0);
      write(32'h00001690, 0);
      write(32'h00001694, 2);
      write(32'h00001698, 5);
      write(32'h0000169C, 4);
      write(32'h000016A0, 11);
      write(32'h000016A4, 16);
      write(32'h000016A8, 14);
      write(32'h000016AC, 6);
      write(32'h000016B0, 11);
      write(32'h000016B4, 10);
      write(32'h000016B8, 1);
      write(32'h000016BC, -5);
      write(32'h000016C0, -6);
      write(32'h000016C4, -6);
      write(32'h000016C8, -6);
      write(32'h000016CC, -3);
      write(32'h000016D0, 2);
      write(32'h000016D4, 11);
      write(32'h000016D8, 16);
      write(32'h000016DC, 12);
      write(32'h000016E0, 6);
      write(32'h000016E4, 10);
      write(32'h000016E8, -1);
      write(32'h000016EC, 0);
      write(32'h000016F0, 0);
      write(32'h000016F4, 0);
      write(32'h000016F8, 0);
      write(32'h000016FC, 0);
      write(32'h00001700, 0);
      write(32'h00001704, 1);
      write(32'h00001708, 4);
      write(32'h0000170C, 4);
      write(32'h00001710, 6);
      write(32'h00001714, 14);
      write(32'h00001718, 12);
      write(32'h0000171C, 13);
      write(32'h00001720, 10);
      write(32'h00001724, 7);
      write(32'h00001728, 3);
      write(32'h0000172C, -4);
      write(32'h00001730, -5);
      write(32'h00001734, -5);
      write(32'h00001738, -5);
      write(32'h0000173C, -5);
      write(32'h00001740, -4);
      write(32'h00001744, 1);
      write(32'h00001748, 5);
      write(32'h0000174C, 2);
      write(32'h00001750, 1);
      write(32'h00001754, 5);
      write(32'h00001758, -1);
      write(32'h0000175C, 0);
      write(32'h00001760, 0);
      write(32'h00001764, 0);
      write(32'h00001768, 0);
      write(32'h0000176C, 0);
      write(32'h00001770, 0);
      write(32'h00001774, 0);
      write(32'h00001778, 3);
      write(32'h0000177C, 6);
      write(32'h00001780, 0);
      write(32'h00001784, 12);
      write(32'h00001788, 14);
      write(32'h0000178C, 11);
      write(32'h00001790, 3);
      write(32'h00001794, 6);
      write(32'h00001798, 2);
      write(32'h0000179C, -5);
      write(32'h000017A0, -4);
      write(32'h000017A4, -5);
      write(32'h000017A8, -6);
      write(32'h000017AC, -8);
      write(32'h000017B0, -9);
      write(32'h000017B4, -10);
      write(32'h000017B8, -4);
      write(32'h000017BC, 0);
      write(32'h000017C0, 1);
      write(32'h000017C4, 2);
      write(32'h000017C8, 0);
      write(32'h000017CC, 0);
      write(32'h000017D0, 0);
      write(32'h000017D4, 0);
      write(32'h000017D8, 0);
      write(32'h000017DC, 0);
      write(32'h000017E0, 0);
      write(32'h000017E4, 0);
      write(32'h000017E8, 3);
      write(32'h000017EC, 8);
      write(32'h000017F0, 0);
      write(32'h000017F4, 8);
      write(32'h000017F8, 14);
      write(32'h000017FC, 8);
      write(32'h00001800, 4);
      write(32'h00001804, 10);
      write(32'h00001808, -1);
      write(32'h0000180C, -6);
      write(32'h00001810, -6);
      write(32'h00001814, -7);
      write(32'h00001818, -9);
      write(32'h0000181C, -12);
      write(32'h00001820, -17);
      write(32'h00001824, -14);
      write(32'h00001828, -5);
      write(32'h0000182C, 4);
      write(32'h00001830, 2);
      write(32'h00001834, 3);
      write(32'h00001838, 0);
      write(32'h0000183C, 0);
      write(32'h00001840, 0);
      write(32'h00001844, 0);
      write(32'h00001848, 0);
      write(32'h0000184C, 0);
      write(32'h00001850, 0);
      write(32'h00001854, -1);
      write(32'h00001858, 1);
      write(32'h0000185C, 9);
      write(32'h00001860, 6);
      write(32'h00001864, 0);
      write(32'h00001868, 9);
      write(32'h0000186C, 6);
      write(32'h00001870, 7);
      write(32'h00001874, 7);
      write(32'h00001878, -1);
      write(32'h0000187C, -4);
      write(32'h00001880, -5);
      write(32'h00001884, -8);
      write(32'h00001888, -10);
      write(32'h0000188C, -18);
      write(32'h00001890, -21);
      write(32'h00001894, -14);
      write(32'h00001898, -5);
      write(32'h0000189C, 6);
      write(32'h000018A0, 5);
      write(32'h000018A4, 5);
      write(32'h000018A8, 2);
      write(32'h000018AC, 0);
      write(32'h000018B0, 0);
      write(32'h000018B4, 0);
      write(32'h000018B8, 0);
      write(32'h000018BC, 0);
      write(32'h000018C0, 0);
      write(32'h000018C4, -1);
      write(32'h000018C8, -1);
      write(32'h000018CC, 8);
      write(32'h000018D0, 10);
      write(32'h000018D4, 3);
      write(32'h000018D8, 0);
      write(32'h000018DC, 1);
      write(32'h000018E0, 6);
      write(32'h000018E4, 5);
      write(32'h000018E8, 1);
      write(32'h000018EC, -4);
      write(32'h000018F0, -5);
      write(32'h000018F4, -8);
      write(32'h000018F8, -14);
      write(32'h000018FC, -18);
      write(32'h00001900, -17);
      write(32'h00001904, -12);
      write(32'h00001908, -2);
      write(32'h0000190C, 5);
      write(32'h00001910, 5);
      write(32'h00001914, 6);
      write(32'h00001918, 3);
      write(32'h0000191C, 0);
      write(32'h00001920, 0);
      write(32'h00001924, 0);
      write(32'h00001928, 0);
      write(32'h0000192C, 0);
      write(32'h00001930, 0);
      write(32'h00001934, -1);
      write(32'h00001938, -3);
      write(32'h0000193C, 6);
      write(32'h00001940, 14);
      write(32'h00001944, 7);
      write(32'h00001948, 0);
      write(32'h0000194C, -2);
      write(32'h00001950, 2);
      write(32'h00001954, 7);
      write(32'h00001958, 0);
      write(32'h0000195C, -5);
      write(32'h00001960, -7);
      write(32'h00001964, -10);
      write(32'h00001968, -15);
      write(32'h0000196C, -13);
      write(32'h00001970, -13);
      write(32'h00001974, -9);
      write(32'h00001978, 0);
      write(32'h0000197C, 4);
      write(32'h00001980, 5);
      write(32'h00001984, 5);
      write(32'h00001988, 1);
      write(32'h0000198C, 0);
      write(32'h00001990, 0);
      write(32'h00001994, 0);
      write(32'h00001998, 0);
      write(32'h0000199C, 0);
      write(32'h000019A0, 0);
      write(32'h000019A4, -1);
      write(32'h000019A8, -2);
      write(32'h000019AC, 0);
      write(32'h000019B0, 14);
      write(32'h000019B4, 18);
      write(32'h000019B8, 11);
      write(32'h000019BC, 2);
      write(32'h000019C0, 7);
      write(32'h000019C4, 13);
      write(32'h000019C8, 4);
      write(32'h000019CC, -4);
      write(32'h000019D0, -6);
      write(32'h000019D4, -7);
      write(32'h000019D8, -11);
      write(32'h000019DC, -12);
      write(32'h000019E0, -12);
      write(32'h000019E4, -7);
      write(32'h000019E8, -3);
      write(32'h000019EC, 2);
      write(32'h000019F0, 5);
      write(32'h000019F4, 1);
      write(32'h000019F8, 0);
      write(32'h000019FC, 0);
      write(32'h00001A00, 0);
      write(32'h00001A04, 0);
      write(32'h00001A08, 0);
      write(32'h00001A0C, 0);
      write(32'h00001A10, 0);
      write(32'h00001A14, 0);
      write(32'h00001A18, -1);
      write(32'h00001A1C, -2);
      write(32'h00001A20, 4);
      write(32'h00001A24, 18);
      write(32'h00001A28, 17);
      write(32'h00001A2C, 11);
      write(32'h00001A30, 14);
      write(32'h00001A34, 13);
      write(32'h00001A38, 5);
      write(32'h00001A3C, -4);
      write(32'h00001A40, -4);
      write(32'h00001A44, -5);
      write(32'h00001A48, -10);
      write(32'h00001A4C, -12);
      write(32'h00001A50, -10);
      write(32'h00001A54, -10);
      write(32'h00001A58, -5);
      write(32'h00001A5C, 0);
      write(32'h00001A60, 1);
      write(32'h00001A64, -1);
      write(32'h00001A68, 0);
      write(32'h00001A6C, 0);
      write(32'h00001A70, 0);
      write(32'h00001A74, 0);
      write(32'h00001A78, 0);
      write(32'h00001A7C, 0);
      write(32'h00001A80, 0);
      write(32'h00001A84, 0);
      write(32'h00001A88, 0);
      write(32'h00001A8C, -2);
      write(32'h00001A90, -3);
      write(32'h00001A94, 5);
      write(32'h00001A98, 16);
      write(32'h00001A9C, 15);
      write(32'h00001AA0, 8);
      write(32'h00001AA4, 7);
      write(32'h00001AA8, -3);
      write(32'h00001AAC, -7);
      write(32'h00001AB0, -7);
      write(32'h00001AB4, -9);
      write(32'h00001AB8, -10);
      write(32'h00001ABC, -11);
      write(32'h00001AC0, -11);
      write(32'h00001AC4, -11);
      write(32'h00001AC8, -7);
      write(32'h00001ACC, -5);
      write(32'h00001AD0, -2);
      write(32'h00001AD4, -1);
      write(32'h00001AD8, 0);
      write(32'h00001ADC, 0);
      write(32'h00001AE0, 0);
      write(32'h00001AE4, 0);
      write(32'h00001AE8, 0);
      write(32'h00001AEC, 0);
      write(32'h00001AF0, 0);
      write(32'h00001AF4, 0);
      write(32'h00001AF8, 0);
      write(32'h00001AFC, -1);
      write(32'h00001B00, -2);
      write(32'h00001B04, -3);
      write(32'h00001B08, 4);
      write(32'h00001B0C, 7);
      write(32'h00001B10, 5);
      write(32'h00001B14, 3);
      write(32'h00001B18, -7);
      write(32'h00001B1C, -8);
      write(32'h00001B20, -9);
      write(32'h00001B24, -10);
      write(32'h00001B28, -11);
      write(32'h00001B2C, -10);
      write(32'h00001B30, -9);
      write(32'h00001B34, -7);
      write(32'h00001B38, -5);
      write(32'h00001B3C, -3);
      write(32'h00001B40, -1);
      write(32'h00001B44, 0);
      write(32'h00001B48, 0);
      write(32'h00001B4C, 0);
      write(32'h00001B50, 0);
      write(32'h00001B54, 0);
      write(32'h00001B58, 0);
      write(32'h00001B5C, 0);
      write(32'h00001B60, 0);
      write(32'h00001B64, 0);
      write(32'h00001B68, 0);
      write(32'h00001B6C, 0);
      write(32'h00001B70, 0);
      write(32'h00001B74, -2);
      write(32'h00001B78, 1);
      write(32'h00001B7C, 8);
      write(32'h00001B80, 8);
      write(32'h00001B84, 5);
      write(32'h00001B88, -4);
      write(32'h00001B8C, -4);
      write(32'h00001B90, -5);
      write(32'h00001B94, -5);
      write(32'h00001B98, -5);
      write(32'h00001B9C, -4);
      write(32'h00001BA0, -4);
      write(32'h00001BA4, -3);
      write(32'h00001BA8, -2);
      write(32'h00001BAC, -1);
      write(32'h00001BB0, 0);
      write(32'h00001BB4, 0);
      write(32'h00001BB8, 0);
      write(32'h00001BBC, 0);
      write(32'h00001BC0, 0);
      write(32'h00001BC4, 0);
      write(32'h00001BC8, 0);
      write(32'h00001BCC, 0);
      write(32'h00001BD0, 0);
      write(32'h00001BD4, 0);
      write(32'h00001BD8, 0);
      write(32'h00001BDC, 0);
      write(32'h00001BE0, 0);
      write(32'h00001BE4, 0);
      write(32'h00001BE8, 0);
      write(32'h00001BEC, 7);
      write(32'h00001BF0, 11);
      write(32'h00001BF4, 7);
      write(32'h00001BF8, -1);
      write(32'h00001BFC, -1);
      write(32'h00001C00, -1);
      write(32'h00001C04, -2);
      write(32'h00001C08, -2);
      write(32'h00001C0C, -2);
      write(32'h00001C10, -2);
      write(32'h00001C14, -1);
      write(32'h00001C18, 0);
      write(32'h00001C1C, 0);
      write(32'h00001C20, 0);
      write(32'h00001C24, 0);
      write(32'h00001C28, 0);
      write(32'h00001C2C, 0);
      write(32'h00001C30, 0);
      write(32'h00001C34, 0);
      write(32'h00001C38, 0);
      write(32'h00001C3C, 0);

      #(PERIOD * 20) ;
      //B
      write(32'h0002E000, -40);
      write(32'h0002E004, 37);
      write(32'h0002E008, 18);
      write(32'h0002E00C, -14);
      write(32'h0002E010, -19);
      write(32'h0002E014, 3);
      write(32'h0002E018, -38);
      write(32'h0002E01C, 43);
      write(32'h0002E020, 20);
      write(32'h0002E024, 56);
      write(32'h0002E028, 0);
      write(32'h0002E02C, 73);
      write(32'h0002E030, -26);
      write(32'h0002E034, 0);
      write(32'h0002E038, -18);
      write(32'h0002E03C, 2);
      write(32'h0002E040, -3);
      write(32'h0002E044, 53);
      write(32'h0002E048, 27);
      write(32'h0002E04C, 15);
      write(32'h0002E050, -15);
      write(32'h0002E054, 21);
      write(32'h0002E058, -29);
      write(32'h0002E05C, -21);
      write(32'h0002E060, 6);
      write(32'h0002E064, -11);
      write(32'h0002E068, 1);
      write(32'h0002E06C, 9);
      write(32'h0002E070, 65);
      write(32'h0002E074, -17);
      write(32'h0002E078, -45);
      write(32'h0002E07C, -9);
      write(32'h0002E080, -23);
      write(32'h0002E084, -20);
      write(32'h0002E088, -25);
      write(32'h0002E08C, 0);
      write(32'h0002E090, -16);
      write(32'h0002E094, 5);
      write(32'h0002E098, 10);
      write(32'h0002E09C, 25);
      write(32'h0002E0A0, -40);
      write(32'h0002E0A4, -12);
      write(32'h0002E0A8, -3);
      write(32'h0002E0AC, -13);
      write(32'h0002E0B0, -37);
      write(32'h0002E0B4, 4);
      #(PERIOD * 20) ;
      //A
      write(32'h00030000, 0);
      write(32'h00030004, 0);
      write(32'h00030008, 0);
      write(32'h0003000C, 0);
      write(32'h00030010, 0);
      write(32'h00030014, 0);
      write(32'h00030018, 0);
      write(32'h0003001C, 0);
      write(32'h00030020, 0);
      write(32'h00030024, 0);
      write(32'h00030028, 0);
      write(32'h0003002C, 0);
      write(32'h00030030, 0);
      write(32'h00030034, 0);
      write(32'h00030038, 0);
      write(32'h0003003C, 0);
      write(32'h00030040, 0);
      write(32'h00030044, 0);
      write(32'h00030048, 0);
      write(32'h0003004C, 0);
      write(32'h00030050, 0);
      write(32'h00030054, 0);
      write(32'h00030058, 0);
      write(32'h0003005C, 0);
      write(32'h00030060, 0);
      write(32'h00030064, 0);
      write(32'h00030068, 0);
      write(32'h0003006C, 0);
      write(32'h00030070, 0);
      write(32'h00030074, 0);
      write(32'h00030078, 0);
      write(32'h0003007C, 0);
      write(32'h00030080, 0);
      write(32'h00030084, 0);
      write(32'h00030088, 0);
      write(32'h0003008C, 0);
      write(32'h00030090, 0);
      write(32'h00030094, 0);
      write(32'h00030098, 0);
      write(32'h0003009C, 0);
      write(32'h000300A0, 0);
      write(32'h000300A4, 0);
      write(32'h000300A8, 0);
      write(32'h000300AC, 0);
      write(32'h000300B0, 0);
      write(32'h000300B4, 0);
      write(32'h000300B8, 0);
      write(32'h000300BC, 0);
      write(32'h000300C0, 0);
      write(32'h000300C4, 0);
      write(32'h000300C8, 0);
      write(32'h000300CC, 0);
      write(32'h000300D0, 0);
      write(32'h000300D4, 0);
      write(32'h000300D8, 0);
      write(32'h000300DC, 0);
      write(32'h000300E0, 0);
      write(32'h000300E4, 0);
      write(32'h000300E8, 0);
      write(32'h000300EC, 0);
      write(32'h000300F0, 0);
      write(32'h000300F4, 0);
      write(32'h000300F8, 0);
      write(32'h000300FC, 0);
      write(32'h00030100, 0);
      write(32'h00030104, 0);
      write(32'h00030108, 0);
      write(32'h0003010C, 0);
      write(32'h00030110, 0);
      write(32'h00030114, 0);
      write(32'h00030118, 0);
      write(32'h0003011C, 0);
      write(32'h00030120, 0);
      write(32'h00030124, 0);
      write(32'h00030128, 0);
      write(32'h0003012C, 0);
      write(32'h00030130, 0);
      write(32'h00030134, 0);
      write(32'h00030138, 0);
      write(32'h0003013C, 0);
      write(32'h00030140, 0);
      write(32'h00030144, 0);
      write(32'h00030148, 0);
      write(32'h0003014C, 0);
      write(32'h00030150, 0);
      write(32'h00030154, 0);
      write(32'h00030158, 0);
      write(32'h0003015C, 0);
      write(32'h00030160, 0);
      write(32'h00030164, 0);
      write(32'h00030168, 0);
      write(32'h0003016C, 0);
      write(32'h00030170, 0);
      write(32'h00030174, 0);
      write(32'h00030178, 0);
      write(32'h0003017C, 0);
      write(32'h00030180, 0);
      write(32'h00030184, 0);
      write(32'h00030188, 0);
      write(32'h0003018C, 0);
      write(32'h00030190, 0);
      write(32'h00030194, 0);
      write(32'h00030198, 0);
      write(32'h0003019C, 0);
      write(32'h000301A0, 0);
      write(32'h000301A4, 0);
      write(32'h000301A8, 0);
      write(32'h000301AC, 0);
      write(32'h000301B0, 0);
      write(32'h000301B4, 0);
      write(32'h000301B8, 0);
      write(32'h000301BC, 0);
      write(32'h000301C0, 0);
      write(32'h000301C4, 0);
      write(32'h000301C8, 0);
      write(32'h000301CC, 0);
      write(32'h000301D0, 0);
      write(32'h000301D4, 0);
      write(32'h000301D8, 0);
      write(32'h000301DC, 0);
      write(32'h000301E0, 0);
      write(32'h000301E4, 0);
      write(32'h000301E8, 0);
      write(32'h000301EC, 0);
      write(32'h000301F0, 0);
      write(32'h000301F4, 0);
      write(32'h000301F8, 0);
      write(32'h000301FC, 0);
      write(32'h00030200, 0);
      write(32'h00030204, 0);
      write(32'h00030208, 0);
      write(32'h0003020C, 0);
      write(32'h00030210, 0);
      write(32'h00030214, 0);
      write(32'h00030218, 0);
      write(32'h0003021C, 0);
      write(32'h00030220, 0);
      write(32'h00030224, 0);
      write(32'h00030228, 0);
      write(32'h0003022C, 0);
      write(32'h00030230, 0);
      write(32'h00030234, 0);
      write(32'h00030238, 0);
      write(32'h0003023C, 0);
      write(32'h00030240, 0);
      write(32'h00030244, 0);
      write(32'h00030248, 0);
      write(32'h0003024C, 0);
      write(32'h00030250, 0);
      write(32'h00030254, 0);
      write(32'h00030258, 0);
      write(32'h0003025C, 0);
      write(32'h00030260, 0);
      write(32'h00030264, 0);
      write(32'h00030268, 0);
      write(32'h0003026C, 0);
      write(32'h00030270, 0);
      write(32'h00030274, 0);
      write(32'h00030278, 0);
      write(32'h0003027C, 0);
      write(32'h00030280, 0);
      write(32'h00030284, 0);
      write(32'h00030288, 0);
      write(32'h0003028C, 0);
      write(32'h00030290, 0);
      write(32'h00030294, 0);
      write(32'h00030298, 0);
      write(32'h0003029C, 0);
      write(32'h000302A0, 0);
      write(32'h000302A4, 0);
      write(32'h000302A8, 0);
      write(32'h000302AC, 0);
      write(32'h000302B0, 0);
      write(32'h000302B4, 0);
      write(32'h000302B8, 0);
      write(32'h000302BC, 0);
      write(32'h000302C0, 0);
      write(32'h000302C4, 0);
      write(32'h000302C8, 0);
      write(32'h000302CC, 0);
      write(32'h000302D0, 0);
      write(32'h000302D4, 0);
      write(32'h000302D8, 0);
      write(32'h000302DC, 0);
      write(32'h000302E0, 0);
      write(32'h000302E4, 0);
      write(32'h000302E8, 0);
      write(32'h000302EC, 0);
      write(32'h000302F0, 0);
      write(32'h000302F4, 0);
      write(32'h000302F8, 0);
      write(32'h000302FC, 0);
      write(32'h00030300, 0);
      write(32'h00030304, 0);
      write(32'h00030308, 0);
      write(32'h0003030C, 0);
      write(32'h00030310, 0);
      write(32'h00030314, 0);
      write(32'h00030318, 0);
      write(32'h0003031C, 0);
      write(32'h00030320, 0);
      write(32'h00030324, 0);
      write(32'h00030328, 0);
      write(32'h0003032C, 0);
      write(32'h00030330, 0);
      write(32'h00030334, 122);
      write(32'h00030338, 169);
      write(32'h0003033C, 79);
      write(32'h00030340, 0);
      write(32'h00030344, 0);
      write(32'h00030348, 0);
      write(32'h0003034C, 0);
      write(32'h00030350, 0);
      write(32'h00030354, 0);
      write(32'h00030358, 0);
      write(32'h0003035C, 0);
      write(32'h00030360, 0);
      write(32'h00030364, 0);
      write(32'h00030368, 0);
      write(32'h0003036C, 0);
      write(32'h00030370, 0);
      write(32'h00030374, 0);
      write(32'h00030378, 0);
      write(32'h0003037C, 0);
      write(32'h00030380, 0);
      write(32'h00030384, 0);
      write(32'h00030388, 0);
      write(32'h0003038C, 0);
      write(32'h00030390, 0);
      write(32'h00030394, 0);
      write(32'h00030398, 0);
      write(32'h0003039C, 0);
      write(32'h000303A0, 0);
      write(32'h000303A4, 197);
      write(32'h000303A8, 255);
      write(32'h000303AC, 115);
      write(32'h000303B0, 0);
      write(32'h000303B4, 0);
      write(32'h000303B8, 0);
      write(32'h000303BC, 0);
      write(32'h000303C0, 0);
      write(32'h000303C4, 0);
      write(32'h000303C8, 0);
      write(32'h000303CC, 0);
      write(32'h000303D0, 0);
      write(32'h000303D4, 0);
      write(32'h000303D8, 0);
      write(32'h000303DC, 0);
      write(32'h000303E0, 0);
      write(32'h000303E4, 0);
      write(32'h000303E8, 0);
      write(32'h000303EC, 0);
      write(32'h000303F0, 0);
      write(32'h000303F4, 0);
      write(32'h000303F8, 0);
      write(32'h000303FC, 0);
      write(32'h00030400, 0);
      write(32'h00030404, 0);
      write(32'h00030408, 0);
      write(32'h0003040C, 0);
      write(32'h00030410, 0);
      write(32'h00030414, 205);
      write(32'h00030418, 255);
      write(32'h0003041C, 116);
      write(32'h00030420, 47);
      write(32'h00030424, 65);
      write(32'h00030428, 92);
      write(32'h0003042C, 124);
      write(32'h00030430, 156);
      write(32'h00030434, 192);
      write(32'h00030438, 134);
      write(32'h0003043C, 0);
      write(32'h00030440, 0);
      write(32'h00030444, 0);
      write(32'h00030448, 0);
      write(32'h0003044C, 0);
      write(32'h00030450, 0);
      write(32'h00030454, 0);
      write(32'h00030458, 0);
      write(32'h0003045C, 0);
      write(32'h00030460, 0);
      write(32'h00030464, 0);
      write(32'h00030468, 0);
      write(32'h0003046C, 0);
      write(32'h00030470, 25);
      write(32'h00030474, 59);
      write(32'h00030478, 90);
      write(32'h0003047C, 121);
      write(32'h00030480, 152);
      write(32'h00030484, 242);
      write(32'h00030488, 255);
      write(32'h0003048C, 239);
      write(32'h00030490, 249);
      write(32'h00030494, 255);
      write(32'h00030498, 255);
      write(32'h0003049C, 255);
      write(32'h000304A0, 255);
      write(32'h000304A4, 250);
      write(32'h000304A8, 186);
      write(32'h000304AC, 0);
      write(32'h000304B0, 0);
      write(32'h000304B4, 0);
      write(32'h000304B8, 0);
      write(32'h000304BC, 0);
      write(32'h000304C0, 0);
      write(32'h000304C4, 0);
      write(32'h000304C8, 0);
      write(32'h000304CC, 0);
      write(32'h000304D0, 0);
      write(32'h000304D4, 0);
      write(32'h000304D8, 0);
      write(32'h000304DC, 0);
      write(32'h000304E0, 171);
      write(32'h000304E4, 255);
      write(32'h000304E8, 255);
      write(32'h000304EC, 255);
      write(32'h000304F0, 255);
      write(32'h000304F4, 255);
      write(32'h000304F8, 255);
      write(32'h000304FC, 228);
      write(32'h00030500, 194);
      write(32'h00030504, 167);
      write(32'h00030508, 141);
      write(32'h0003050C, 111);
      write(32'h00030510, 80);
      write(32'h00030514, 50);
      write(32'h00030518, 19);
      write(32'h0003051C, 0);
      write(32'h00030520, 0);
      write(32'h00030524, 0);
      write(32'h00030528, 0);
      write(32'h0003052C, 0);
      write(32'h00030530, 0);
      write(32'h00030534, 0);
      write(32'h00030538, 0);
      write(32'h0003053C, 0);
      write(32'h00030540, 0);
      write(32'h00030544, 0);
      write(32'h00030548, 0);
      write(32'h0003054C, 0);
      write(32'h00030550, 107);
      write(32'h00030554, 174);
      write(32'h00030558, 137);
      write(32'h0003055C, 103);
      write(32'h00030560, 71);
      write(32'h00030564, 228);
      write(32'h00030568, 253);
      write(32'h0003056C, 84);
      write(32'h00030570, 9);
      write(32'h00030574, 0);
      write(32'h00030578, 0);
      write(32'h0003057C, 0);
      write(32'h00030580, 0);
      write(32'h00030584, 0);
      write(32'h00030588, 0);
      write(32'h0003058C, 0);
      write(32'h00030590, 0);
      write(32'h00030594, 0);
      write(32'h00030598, 0);
      write(32'h0003059C, 0);
      write(32'h000305A0, 0);
      write(32'h000305A4, 0);
      write(32'h000305A8, 0);
      write(32'h000305AC, 0);
      write(32'h000305B0, 0);
      write(32'h000305B4, 0);
      write(32'h000305B8, 0);
      write(32'h000305BC, 0);
      write(32'h000305C0, 0);
      write(32'h000305C4, 0);
      write(32'h000305C8, 0);
      write(32'h000305CC, 0);
      write(32'h000305D0, 0);
      write(32'h000305D4, 218);
      write(32'h000305D8, 255);
      write(32'h000305DC, 81);
      write(32'h000305E0, 12);
      write(32'h000305E4, 13);
      write(32'h000305E8, 13);
      write(32'h000305EC, 8);
      write(32'h000305F0, 0);
      write(32'h000305F4, 0);
      write(32'h000305F8, 0);
      write(32'h000305FC, 0);
      write(32'h00030600, 0);
      write(32'h00030604, 0);
      write(32'h00030608, 0);
      write(32'h0003060C, 0);
      write(32'h00030610, 0);
      write(32'h00030614, 0);
      write(32'h00030618, 0);
      write(32'h0003061C, 0);
      write(32'h00030620, 0);
      write(32'h00030624, 0);
      write(32'h00030628, 0);
      write(32'h0003062C, 0);
      write(32'h00030630, 0);
      write(32'h00030634, 0);
      write(32'h00030638, 0);
      write(32'h0003063C, 10);
      write(32'h00030640, 80);
      write(32'h00030644, 234);
      write(32'h00030648, 255);
      write(32'h0003064C, 250);
      write(32'h00030650, 247);
      write(32'h00030654, 247);
      write(32'h00030658, 232);
      write(32'h0003065C, 203);
      write(32'h00030660, 145);
      write(32'h00030664, 64);
      write(32'h00030668, 0);
      write(32'h0003066C, 0);
      write(32'h00030670, 0);
      write(32'h00030674, 0);
      write(32'h00030678, 0);
      write(32'h0003067C, 0);
      write(32'h00030680, 0);
      write(32'h00030684, 0);
      write(32'h00030688, 0);
      write(32'h0003068C, 0);
      write(32'h00030690, 0);
      write(32'h00030694, 0);
      write(32'h00030698, 0);
      write(32'h0003069C, 0);
      write(32'h000306A0, 0);
      write(32'h000306A4, 0);
      write(32'h000306A8, 76);
      write(32'h000306AC, 200);
      write(32'h000306B0, 255);
      write(32'h000306B4, 255);
      write(32'h000306B8, 254);
      write(32'h000306BC, 225);
      write(32'h000306C0, 211);
      write(32'h000306C4, 211);
      write(32'h000306C8, 251);
      write(32'h000306CC, 255);
      write(32'h000306D0, 255);
      write(32'h000306D4, 250);
      write(32'h000306D8, 156);
      write(32'h000306DC, 21);
      write(32'h000306E0, 0);
      write(32'h000306E4, 0);
      write(32'h000306E8, 0);
      write(32'h000306EC, 0);
      write(32'h000306F0, 0);
      write(32'h000306F4, 0);
      write(32'h000306F8, 0);
      write(32'h000306FC, 0);
      write(32'h00030700, 0);
      write(32'h00030704, 0);
      write(32'h00030708, 0);
      write(32'h0003070C, 0);
      write(32'h00030710, 3);
      write(32'h00030714, 124);
      write(32'h00030718, 251);
      write(32'h0003071C, 255);
      write(32'h00030720, 155);
      write(32'h00030724, 230);
      write(32'h00030728, 253);
      write(32'h0003072C, 82);
      write(32'h00030730, 0);
      write(32'h00030734, 27);
      write(32'h00030738, 238);
      write(32'h0003073C, 251);
      write(32'h00030740, 144);
      write(32'h00030744, 200);
      write(32'h00030748, 255);
      write(32'h0003074C, 193);
      write(32'h00030750, 22);
      write(32'h00030754, 0);
      write(32'h00030758, 0);
      write(32'h0003075C, 0);
      write(32'h00030760, 0);
      write(32'h00030764, 0);
      write(32'h00030768, 0);
      write(32'h0003076C, 0);
      write(32'h00030770, 0);
      write(32'h00030774, 0);
      write(32'h00030778, 0);
      write(32'h0003077C, 0);
      write(32'h00030780, 118);
      write(32'h00030784, 255);
      write(32'h00030788, 239);
      write(32'h0003078C, 86);
      write(32'h00030790, 0);
      write(32'h00030794, 202);
      write(32'h00030798, 255);
      write(32'h0003079C, 102);
      write(32'h000307A0, 0);
      write(32'h000307A4, 115);
      write(32'h000307A8, 255);
      write(32'h000307AC, 217);
      write(32'h000307B0, 10);
      write(32'h000307B4, 24);
      write(32'h000307B8, 198);
      write(32'h000307BC, 255);
      write(32'h000307C0, 147);
      write(32'h000307C4, 1);
      write(32'h000307C8, 0);
      write(32'h000307CC, 0);
      write(32'h000307D0, 0);
      write(32'h000307D4, 0);
      write(32'h000307D8, 0);
      write(32'h000307DC, 0);
      write(32'h000307E0, 0);
      write(32'h000307E4, 0);
      write(32'h000307E8, 0);
      write(32'h000307EC, 54);
      write(32'h000307F0, 242);
      write(32'h000307F4, 251);
      write(32'h000307F8, 90);
      write(32'h000307FC, 0);
      write(32'h00030800, 0);
      write(32'h00030804, 185);
      write(32'h00030808, 255);
      write(32'h0003080C, 115);
      write(32'h00030810, 8);
      write(32'h00030814, 204);
      write(32'h00030818, 255);
      write(32'h0003081C, 126);
      write(32'h00030820, 0);
      write(32'h00030824, 0);
      write(32'h00030828, 65);
      write(32'h0003082C, 252);
      write(32'h00030830, 230);
      write(32'h00030834, 35);
      write(32'h00030838, 0);
      write(32'h0003083C, 0);
      write(32'h00030840, 0);
      write(32'h00030844, 0);
      write(32'h00030848, 0);
      write(32'h0003084C, 0);
      write(32'h00030850, 0);
      write(32'h00030854, 0);
      write(32'h00030858, 0);
      write(32'h0003085C, 149);
      write(32'h00030860, 255);
      write(32'h00030864, 167);
      write(32'h00030868, 2);
      write(32'h0003086C, 0);
      write(32'h00030870, 0);
      write(32'h00030874, 163);
      write(32'h00030878, 255);
      write(32'h0003087C, 129);
      write(32'h00030880, 83);
      write(32'h00030884, 255);
      write(32'h00030888, 229);
      write(32'h0003088C, 30);
      write(32'h00030890, 0);
      write(32'h00030894, 0);
      write(32'h00030898, 17);
      write(32'h0003089C, 214);
      write(32'h000308A0, 255);
      write(32'h000308A4, 67);
      write(32'h000308A8, 0);
      write(32'h000308AC, 0);
      write(32'h000308B0, 0);
      write(32'h000308B4, 0);
      write(32'h000308B8, 0);
      write(32'h000308BC, 0);
      write(32'h000308C0, 0);
      write(32'h000308C4, 0);
      write(32'h000308C8, 5);
      write(32'h000308CC, 212);
      write(32'h000308D0, 254);
      write(32'h000308D4, 88);
      write(32'h000308D8, 0);
      write(32'h000308DC, 0);
      write(32'h000308E0, 0);
      write(32'h000308E4, 137);
      write(32'h000308E8, 255);
      write(32'h000308EC, 188);
      write(32'h000308F0, 214);
      write(32'h000308F4, 255);
      write(32'h000308F8, 112);
      write(32'h000308FC, 0);
      write(32'h00030900, 0);
      write(32'h00030904, 0);
      write(32'h00030908, 14);
      write(32'h0003090C, 203);
      write(32'h00030910, 255);
      write(32'h00030914, 71);
      write(32'h00030918, 0);
      write(32'h0003091C, 0);
      write(32'h00030920, 0);
      write(32'h00030924, 0);
      write(32'h00030928, 0);
      write(32'h0003092C, 0);
      write(32'h00030930, 0);
      write(32'h00030934, 0);
      write(32'h00030938, 7);
      write(32'h0003093C, 232);
      write(32'h00030940, 249);
      write(32'h00030944, 63);
      write(32'h00030948, 0);
      write(32'h0003094C, 0);
      write(32'h00030950, 0);
      write(32'h00030954, 105);
      write(32'h00030958, 255);
      write(32'h0003095C, 255);
      write(32'h00030960, 255);
      write(32'h00030964, 173);
      write(32'h00030968, 7);
      write(32'h0003096C, 0);
      write(32'h00030970, 0);
      write(32'h00030974, 0);
      write(32'h00030978, 38);
      write(32'h0003097C, 244);
      write(32'h00030980, 239);
      write(32'h00030984, 46);
      write(32'h00030988, 0);
      write(32'h0003098C, 0);
      write(32'h00030990, 0);
      write(32'h00030994, 0);
      write(32'h00030998, 0);
      write(32'h0003099C, 0);
      write(32'h000309A0, 0);
      write(32'h000309A4, 0);
      write(32'h000309A8, 4);
      write(32'h000309AC, 207);
      write(32'h000309B0, 255);
      write(32'h000309B4, 107);
      write(32'h000309B8, 0);
      write(32'h000309BC, 0);
      write(32'h000309C0, 0);
      write(32'h000309C4, 106);
      write(32'h000309C8, 255);
      write(32'h000309CC, 255);
      write(32'h000309D0, 187);
      write(32'h000309D4, 25);
      write(32'h000309D8, 0);
      write(32'h000309DC, 0);
      write(32'h000309E0, 0);
      write(32'h000309E4, 0);
      write(32'h000309E8, 152);
      write(32'h000309EC, 255);
      write(32'h000309F0, 182);
      write(32'h000309F4, 7);
      write(32'h000309F8, 0);
      write(32'h000309FC, 0);
      write(32'h00030A00, 0);
      write(32'h00030A04, 0);
      write(32'h00030A08, 0);
      write(32'h00030A0C, 0);
      write(32'h00030A10, 0);
      write(32'h00030A14, 0);
      write(32'h00030A18, 0);
      write(32'h00030A1C, 119);
      write(32'h00030A20, 255);
      write(32'h00030A24, 231);
      write(32'h00030A28, 103);
      write(32'h00030A2C, 75);
      write(32'h00030A30, 155);
      write(32'h00030A34, 243);
      write(32'h00030A38, 255);
      write(32'h00030A3C, 255);
      write(32'h00030A40, 105);
      write(32'h00030A44, 0);
      write(32'h00030A48, 0);
      write(32'h00030A4C, 0);
      write(32'h00030A50, 5);
      write(32'h00030A54, 125);
      write(32'h00030A58, 253);
      write(32'h00030A5C, 244);
      write(32'h00030A60, 62);
      write(32'h00030A64, 0);
      write(32'h00030A68, 0);
      write(32'h00030A6C, 0);
      write(32'h00030A70, 0);
      write(32'h00030A74, 0);
      write(32'h00030A78, 0);
      write(32'h00030A7C, 0);
      write(32'h00030A80, 0);
      write(32'h00030A84, 0);
      write(32'h00030A88, 0);
      write(32'h00030A8C, 15);
      write(32'h00030A90, 167);
      write(32'h00030A94, 254);
      write(32'h00030A98, 255);
      write(32'h00030A9C, 255);
      write(32'h00030AA0, 255);
      write(32'h00030AA4, 212);
      write(32'h00030AA8, 211);
      write(32'h00030AAC, 247);
      write(32'h00030AB0, 131);
      write(32'h00030AB4, 0);
      write(32'h00030AB8, 0);
      write(32'h00030ABC, 41);
      write(32'h00030AC0, 168);
      write(32'h00030AC4, 255);
      write(32'h00030AC8, 250);
      write(32'h00030ACC, 105);
      write(32'h00030AD0, 0);
      write(32'h00030AD4, 0);
      write(32'h00030AD8, 0);
      write(32'h00030ADC, 0);
      write(32'h00030AE0, 0);
      write(32'h00030AE4, 0);
      write(32'h00030AE8, 0);
      write(32'h00030AEC, 0);
      write(32'h00030AF0, 0);
      write(32'h00030AF4, 0);
      write(32'h00030AF8, 0);
      write(32'h00030AFC, 0);
      write(32'h00030B00, 5);
      write(32'h00030B04, 83);
      write(32'h00030B08, 138);
      write(32'h00030B0C, 136);
      write(32'h00030B10, 91);
      write(32'h00030B14, 14);
      write(32'h00030B18, 59);
      write(32'h00030B1C, 64);
      write(32'h00030B20, 5);
      write(32'h00030B24, 3);
      write(32'h00030B28, 119);
      write(32'h00030B2C, 236);
      write(32'h00030B30, 255);
      write(32'h00030B34, 241);
      write(32'h00030B38, 103);
      write(32'h00030B3C, 0);
      write(32'h00030B40, 0);
      write(32'h00030B44, 0);
      write(32'h00030B48, 0);
      write(32'h00030B4C, 0);
      write(32'h00030B50, 0);
      write(32'h00030B54, 0);
      write(32'h00030B58, 0);
      write(32'h00030B5C, 0);
      write(32'h00030B60, 0);
      write(32'h00030B64, 0);
      write(32'h00030B68, 0);
      write(32'h00030B6C, 0);
      write(32'h00030B70, 0);
      write(32'h00030B74, 0);
      write(32'h00030B78, 0);
      write(32'h00030B7C, 0);
      write(32'h00030B80, 0);
      write(32'h00030B84, 0);
      write(32'h00030B88, 0);
      write(32'h00030B8C, 0);
      write(32'h00030B90, 0);
      write(32'h00030B94, 2);
      write(32'h00030B98, 116);
      write(32'h00030B9C, 242);
      write(32'h00030BA0, 186);
      write(32'h00030BA4, 58);
      write(32'h00030BA8, 0);
      write(32'h00030BAC, 0);
      write(32'h00030BB0, 0);
      write(32'h00030BB4, 0);
      write(32'h00030BB8, 0);
      write(32'h00030BBC, 0);
      write(32'h00030BC0, 0);
      write(32'h00030BC4, 0);
      write(32'h00030BC8, 0);
      write(32'h00030BCC, 0);
      write(32'h00030BD0, 0);
      write(32'h00030BD4, 0);
      write(32'h00030BD8, 0);
      write(32'h00030BDC, 0);
      write(32'h00030BE0, 0);
      write(32'h00030BE4, 0);
      write(32'h00030BE8, 0);
      write(32'h00030BEC, 0);
      write(32'h00030BF0, 0);
      write(32'h00030BF4, 0);
      write(32'h00030BF8, 0);
      write(32'h00030BFC, 0);
      write(32'h00030C00, 0);
      write(32'h00030C04, 0);
      write(32'h00030C08, 6);
      write(32'h00030C0C, 62);
      write(32'h00030C10, 7);
      write(32'h00030C14, 0);
      write(32'h00030C18, 0);
      write(32'h00030C1C, 0);
      write(32'h00030C20, 0);
      write(32'h00030C24, 0);
      write(32'h00030C28, 0);
      write(32'h00030C2C, 0);
      write(32'h00030C30, 0);
      write(32'h00030C34, 0);
      write(32'h00030C38, 0);
      write(32'h00030C3C, 0);

      $display("DATA A");

      #(PERIOD * 200) ;
      
      //I
      write(32'h00030000, 0);
      write(32'h00030004, 0);
      write(32'h00030008, 0);
      write(32'h0003000C, 0);
      write(32'h00030010, 0);
      write(32'h00030014, 0);
      write(32'h00030018, 0);
      write(32'h0003001C, 0);
      write(32'h00030020, 0);
      write(32'h00030024, 0);
      write(32'h00030028, 0);
      write(32'h0003002C, 0);
      write(32'h00030030, 0);
      write(32'h00030034, 0);
      write(32'h00030038, 0);
      write(32'h0003003C, 0);
      write(32'h00030040, 0);
      write(32'h00030044, 0);
      write(32'h00030048, 0);
      write(32'h0003004C, 0);
      write(32'h00030050, 0);
      write(32'h00030054, 0);
      write(32'h00030058, 0);
      write(32'h0003005C, 0);
      write(32'h00030060, 0);
      write(32'h00030064, 0);
      write(32'h00030068, 0);
      write(32'h0003006C, 0);
      write(32'h00030070, 0);
      write(32'h00030074, 0);
      write(32'h00030078, 0);
      write(32'h0003007C, 0);
      write(32'h00030080, 0);
      write(32'h00030084, 0);
      write(32'h00030088, 0);
      write(32'h0003008C, 0);
      write(32'h00030090, 0);
      write(32'h00030094, 0);
      write(32'h00030098, 0);
      write(32'h0003009C, 0);
      write(32'h000300A0, 0);
      write(32'h000300A4, 0);
      write(32'h000300A8, 0);
      write(32'h000300AC, 0);
      write(32'h000300B0, 0);
      write(32'h000300B4, 0);
      write(32'h000300B8, 0);
      write(32'h000300BC, 0);
      write(32'h000300C0, 0);
      write(32'h000300C4, 0);
      write(32'h000300C8, 0);
      write(32'h000300CC, 0);
      write(32'h000300D0, 0);
      write(32'h000300D4, 0);
      write(32'h000300D8, 0);
      write(32'h000300DC, 0);
      write(32'h000300E0, 0);
      write(32'h000300E4, 0);
      write(32'h000300E8, 0);
      write(32'h000300EC, 0);
      write(32'h000300F0, 0);
      write(32'h000300F4, 0);
      write(32'h000300F8, 0);
      write(32'h000300FC, 0);
      write(32'h00030100, 0);
      write(32'h00030104, 0);
      write(32'h00030108, 0);
      write(32'h0003010C, 0);
      write(32'h00030110, 0);
      write(32'h00030114, 0);
      write(32'h00030118, 0);
      write(32'h0003011C, 0);
      write(32'h00030120, 0);
      write(32'h00030124, 0);
      write(32'h00030128, 0);
      write(32'h0003012C, 0);
      write(32'h00030130, 0);
      write(32'h00030134, 0);
      write(32'h00030138, 0);
      write(32'h0003013C, 0);
      write(32'h00030140, 0);
      write(32'h00030144, 0);
      write(32'h00030148, 0);
      write(32'h0003014C, 0);
      write(32'h00030150, 0);
      write(32'h00030154, 0);
      write(32'h00030158, 0);
      write(32'h0003015C, 0);
      write(32'h00030160, 0);
      write(32'h00030164, 0);
      write(32'h00030168, 0);
      write(32'h0003016C, 0);
      write(32'h00030170, 0);
      write(32'h00030174, 0);
      write(32'h00030178, 0);
      write(32'h0003017C, 0);
      write(32'h00030180, 0);
      write(32'h00030184, 0);
      write(32'h00030188, 0);
      write(32'h0003018C, 0);
      write(32'h00030190, 0);
      write(32'h00030194, 0);
      write(32'h00030198, 0);
      write(32'h0003019C, 0);
      write(32'h000301A0, 0);
      write(32'h000301A4, 0);
      write(32'h000301A8, 0);
      write(32'h000301AC, 0);
      write(32'h000301B0, 0);
      write(32'h000301B4, 0);
      write(32'h000301B8, 0);
      write(32'h000301BC, 0);
      write(32'h000301C0, 0);
      write(32'h000301C4, 0);
      write(32'h000301C8, 0);
      write(32'h000301CC, 0);
      write(32'h000301D0, 0);
      write(32'h000301D4, 0);
      write(32'h000301D8, 0);
      write(32'h000301DC, 0);
      write(32'h000301E0, 0);
      write(32'h000301E4, 0);
      write(32'h000301E8, 0);
      write(32'h000301EC, 0);
      write(32'h000301F0, 0);
      write(32'h000301F4, 0);
      write(32'h000301F8, 0);
      write(32'h000301FC, 0);
      write(32'h00030200, 0);
      write(32'h00030204, 0);
      write(32'h00030208, 0);
      write(32'h0003020C, 0);
      write(32'h00030210, 0);
      write(32'h00030214, 0);
      write(32'h00030218, 0);
      write(32'h0003021C, 0);
      write(32'h00030220, 0);
      write(32'h00030224, 0);
      write(32'h00030228, 0);
      write(32'h0003022C, 0);
      write(32'h00030230, 0);
      write(32'h00030234, 0);
      write(32'h00030238, 0);
      write(32'h0003023C, 0);
      write(32'h00030240, 0);
      write(32'h00030244, 0);
      write(32'h00030248, 0);
      write(32'h0003024C, 0);
      write(32'h00030250, 0);
      write(32'h00030254, 0);
      write(32'h00030258, 0);
      write(32'h0003025C, 0);
      write(32'h00030260, 0);
      write(32'h00030264, 0);
      write(32'h00030268, 0);
      write(32'h0003026C, 0);
      write(32'h00030270, 0);
      write(32'h00030274, 0);
      write(32'h00030278, 0);
      write(32'h0003027C, 0);
      write(32'h00030280, 0);
      write(32'h00030284, 0);
      write(32'h00030288, 0);
      write(32'h0003028C, 0);
      write(32'h00030290, 0);
      write(32'h00030294, 0);
      write(32'h00030298, 0);
      write(32'h0003029C, 0);
      write(32'h000302A0, 0);
      write(32'h000302A4, 0);
      write(32'h000302A8, 0);
      write(32'h000302AC, 0);
      write(32'h000302B0, 0);
      write(32'h000302B4, 0);
      write(32'h000302B8, 0);
      write(32'h000302BC, 0);
      write(32'h000302C0, 0);
      write(32'h000302C4, 0);
      write(32'h000302C8, 0);
      write(32'h000302CC, 0);
      write(32'h000302D0, 0);
      write(32'h000302D4, 0);
      write(32'h000302D8, 0);
      write(32'h000302DC, 0);
      write(32'h000302E0, 0);
      write(32'h000302E4, 0);
      write(32'h000302E8, 0);
      write(32'h000302EC, 0);
      write(32'h000302F0, 0);
      write(32'h000302F4, 0);
      write(32'h000302F8, 0);
      write(32'h000302FC, 0);
      write(32'h00030300, 0);
      write(32'h00030304, 0);
      write(32'h00030308, 0);
      write(32'h0003030C, 0);
      write(32'h00030310, 0);
      write(32'h00030314, 0);
      write(32'h00030318, 0);
      write(32'h0003031C, 5);
      write(32'h00030320, 17);
      write(32'h00030324, 4);
      write(32'h00030328, 0);
      write(32'h0003032C, 0);
      write(32'h00030330, 0);
      write(32'h00030334, 0);
      write(32'h00030338, 0);
      write(32'h0003033C, 0);
      write(32'h00030340, 0);
      write(32'h00030344, 0);
      write(32'h00030348, 0);
      write(32'h0003034C, 0);
      write(32'h00030350, 0);
      write(32'h00030354, 0);
      write(32'h00030358, 0);
      write(32'h0003035C, 0);
      write(32'h00030360, 0);
      write(32'h00030364, 0);
      write(32'h00030368, 0);
      write(32'h0003036C, 0);
      write(32'h00030370, 0);
      write(32'h00030374, 0);
      write(32'h00030378, 0);
      write(32'h0003037C, 0);
      write(32'h00030380, 0);
      write(32'h00030384, 0);
      write(32'h00030388, 0);
      write(32'h0003038C, 46);
      write(32'h00030390, 205);
      write(32'h00030394, 167);
      write(32'h00030398, 15);
      write(32'h0003039C, 0);
      write(32'h000303A0, 0);
      write(32'h000303A4, 0);
      write(32'h000303A8, 0);
      write(32'h000303AC, 0);
      write(32'h000303B0, 0);
      write(32'h000303B4, 0);
      write(32'h000303B8, 0);
      write(32'h000303BC, 1);
      write(32'h000303C0, 53);
      write(32'h000303C4, 53);
      write(32'h000303C8, 0);
      write(32'h000303CC, 0);
      write(32'h000303D0, 0);
      write(32'h000303D4, 0);
      write(32'h000303D8, 0);
      write(32'h000303DC, 0);
      write(32'h000303E0, 0);
      write(32'h000303E4, 0);
      write(32'h000303E8, 0);
      write(32'h000303EC, 0);
      write(32'h000303F0, 0);
      write(32'h000303F4, 0);
      write(32'h000303F8, 0);
      write(32'h000303FC, 60);
      write(32'h00030400, 252);
      write(32'h00030404, 239);
      write(32'h00030408, 23);
      write(32'h0003040C, 0);
      write(32'h00030410, 0);
      write(32'h00030414, 0);
      write(32'h00030418, 0);
      write(32'h0003041C, 0);
      write(32'h00030420, 0);
      write(32'h00030424, 0);
      write(32'h00030428, 0);
      write(32'h0003042C, 124);
      write(32'h00030430, 240);
      write(32'h00030434, 190);
      write(32'h00030438, 8);
      write(32'h0003043C, 0);
      write(32'h00030440, 0);
      write(32'h00030444, 0);
      write(32'h00030448, 0);
      write(32'h0003044C, 0);
      write(32'h00030450, 0);
      write(32'h00030454, 0);
      write(32'h00030458, 0);
      write(32'h0003045C, 0);
      write(32'h00030460, 0);
      write(32'h00030464, 0);
      write(32'h00030468, 0);
      write(32'h0003046C, 72);
      write(32'h00030470, 255);
      write(32'h00030474, 212);
      write(32'h00030478, 16);
      write(32'h0003047C, 0);
      write(32'h00030480, 0);
      write(32'h00030484, 0);
      write(32'h00030488, 0);
      write(32'h0003048C, 0);
      write(32'h00030490, 0);
      write(32'h00030494, 0);
      write(32'h00030498, 0);
      write(32'h0003049C, 69);
      write(32'h000304A0, 252);
      write(32'h000304A4, 249);
      write(32'h000304A8, 65);
      write(32'h000304AC, 0);
      write(32'h000304B0, 0);
      write(32'h000304B4, 0);
      write(32'h000304B8, 0);
      write(32'h000304BC, 0);
      write(32'h000304C0, 0);
      write(32'h000304C4, 0);
      write(32'h000304C8, 0);
      write(32'h000304CC, 0);
      write(32'h000304D0, 0);
      write(32'h000304D4, 0);
      write(32'h000304D8, 0);
      write(32'h000304DC, 78);
      write(32'h000304E0, 255);
      write(32'h000304E4, 199);
      write(32'h000304E8, 13);
      write(32'h000304EC, 0);
      write(32'h000304F0, 0);
      write(32'h000304F4, 0);
      write(32'h000304F8, 0);
      write(32'h000304FC, 0);
      write(32'h00030500, 0);
      write(32'h00030504, 0);
      write(32'h00030508, 0);
      write(32'h0003050C, 6);
      write(32'h00030510, 178);
      write(32'h00030514, 255);
      write(32'h00030518, 157);
      write(32'h0003051C, 0);
      write(32'h00030520, 0);
      write(32'h00030524, 0);
      write(32'h00030528, 0);
      write(32'h0003052C, 0);
      write(32'h00030530, 0);
      write(32'h00030534, 0);
      write(32'h00030538, 0);
      write(32'h0003053C, 0);
      write(32'h00030540, 0);
      write(32'h00030544, 0);
      write(32'h00030548, 0);
      write(32'h0003054C, 83);
      write(32'h00030550, 255);
      write(32'h00030554, 191);
      write(32'h00030558, 10);
      write(32'h0003055C, 0);
      write(32'h00030560, 0);
      write(32'h00030564, 0);
      write(32'h00030568, 0);
      write(32'h0003056C, 0);
      write(32'h00030570, 0);
      write(32'h00030574, 0);
      write(32'h00030578, 0);
      write(32'h0003057C, 0);
      write(32'h00030580, 78);
      write(32'h00030584, 254);
      write(32'h00030588, 230);
      write(32'h0003058C, 27);
      write(32'h00030590, 0);
      write(32'h00030594, 0);
      write(32'h00030598, 0);
      write(32'h0003059C, 0);
      write(32'h000305A0, 0);
      write(32'h000305A4, 0);
      write(32'h000305A8, 0);
      write(32'h000305AC, 0);
      write(32'h000305B0, 0);
      write(32'h000305B4, 0);
      write(32'h000305B8, 0);
      write(32'h000305BC, 85);
      write(32'h000305C0, 255);
      write(32'h000305C4, 188);
      write(32'h000305C8, 9);
      write(32'h000305CC, 0);
      write(32'h000305D0, 0);
      write(32'h000305D4, 0);
      write(32'h000305D8, 0);
      write(32'h000305DC, 0);
      write(32'h000305E0, 0);
      write(32'h000305E4, 0);
      write(32'h000305E8, 0);
      write(32'h000305EC, 0);
      write(32'h000305F0, 8);
      write(32'h000305F4, 209);
      write(32'h000305F8, 254);
      write(32'h000305FC, 98);
      write(32'h00030600, 0);
      write(32'h00030604, 0);
      write(32'h00030608, 0);
      write(32'h0003060C, 0);
      write(32'h00030610, 0);
      write(32'h00030614, 0);
      write(32'h00030618, 0);
      write(32'h0003061C, 0);
      write(32'h00030620, 0);
      write(32'h00030624, 0);
      write(32'h00030628, 0);
      write(32'h0003062C, 80);
      write(32'h00030630, 255);
      write(32'h00030634, 191);
      write(32'h00030638, 10);
      write(32'h0003063C, 0);
      write(32'h00030640, 0);
      write(32'h00030644, 0);
      write(32'h00030648, 0);
      write(32'h0003064C, 0);
      write(32'h00030650, 0);
      write(32'h00030654, 0);
      write(32'h00030658, 0);
      write(32'h0003065C, 0);
      write(32'h00030660, 0);
      write(32'h00030664, 125);
      write(32'h00030668, 255);
      write(32'h0003066C, 167);
      write(32'h00030670, 3);
      write(32'h00030674, 0);
      write(32'h00030678, 0);
      write(32'h0003067C, 0);
      write(32'h00030680, 0);
      write(32'h00030684, 0);
      write(32'h00030688, 0);
      write(32'h0003068C, 0);
      write(32'h00030690, 0);
      write(32'h00030694, 0);
      write(32'h00030698, 0);
      write(32'h0003069C, 73);
      write(32'h000306A0, 255);
      write(32'h000306A4, 202);
      write(32'h000306A8, 13);
      write(32'h000306AC, 0);
      write(32'h000306B0, 0);
      write(32'h000306B4, 0);
      write(32'h000306B8, 0);
      write(32'h000306BC, 0);
      write(32'h000306C0, 0);
      write(32'h000306C4, 0);
      write(32'h000306C8, 0);
      write(32'h000306CC, 0);
      write(32'h000306D0, 0);
      write(32'h000306D4, 59);
      write(32'h000306D8, 246);
      write(32'h000306DC, 232);
      write(32'h000306E0, 23);
      write(32'h000306E4, 0);
      write(32'h000306E8, 0);
      write(32'h000306EC, 0);
      write(32'h000306F0, 0);
      write(32'h000306F4, 0);
      write(32'h000306F8, 0);
      write(32'h000306FC, 0);
      write(32'h00030700, 0);
      write(32'h00030704, 0);
      write(32'h00030708, 0);
      write(32'h0003070C, 58);
      write(32'h00030710, 248);
      write(32'h00030714, 223);
      write(32'h00030718, 19);
      write(32'h0003071C, 0);
      write(32'h00030720, 0);
      write(32'h00030724, 0);
      write(32'h00030728, 0);
      write(32'h0003072C, 0);
      write(32'h00030730, 0);
      write(32'h00030734, 0);
      write(32'h00030738, 0);
      write(32'h0003073C, 0);
      write(32'h00030740, 0);
      write(32'h00030744, 15);
      write(32'h00030748, 211);
      write(32'h0003074C, 255);
      write(32'h00030750, 68);
      write(32'h00030754, 0);
      write(32'h00030758, 0);
      write(32'h0003075C, 0);
      write(32'h00030760, 0);
      write(32'h00030764, 0);
      write(32'h00030768, 0);
      write(32'h0003076C, 0);
      write(32'h00030770, 0);
      write(32'h00030774, 0);
      write(32'h00030778, 0);
      write(32'h0003077C, 36);
      write(32'h00030780, 229);
      write(32'h00030784, 249);
      write(32'h00030788, 30);
      write(32'h0003078C, 0);
      write(32'h00030790, 0);
      write(32'h00030794, 0);
      write(32'h00030798, 0);
      write(32'h0003079C, 0);
      write(32'h000307A0, 0);
      write(32'h000307A4, 0);
      write(32'h000307A8, 0);
      write(32'h000307AC, 0);
      write(32'h000307B0, 0);
      write(32'h000307B4, 0);
      write(32'h000307B8, 171);
      write(32'h000307BC, 255);
      write(32'h000307C0, 125);
      write(32'h000307C4, 0);
      write(32'h000307C8, 0);
      write(32'h000307CC, 0);
      write(32'h000307D0, 0);
      write(32'h000307D4, 0);
      write(32'h000307D8, 0);
      write(32'h000307DC, 0);
      write(32'h000307E0, 0);
      write(32'h000307E4, 0);
      write(32'h000307E8, 0);
      write(32'h000307EC, 11);
      write(32'h000307F0, 206);
      write(32'h000307F4, 255);
      write(32'h000307F8, 67);
      write(32'h000307FC, 0);
      write(32'h00030800, 0);
      write(32'h00030804, 0);
      write(32'h00030808, 0);
      write(32'h0003080C, 0);
      write(32'h00030810, 0);
      write(32'h00030814, 0);
      write(32'h00030818, 0);
      write(32'h0003081C, 0);
      write(32'h00030820, 0);
      write(32'h00030824, 0);
      write(32'h00030828, 121);
      write(32'h0003082C, 255);
      write(32'h00030830, 172);
      write(32'h00030834, 0);
      write(32'h00030838, 0);
      write(32'h0003083C, 0);
      write(32'h00030840, 0);
      write(32'h00030844, 0);
      write(32'h00030848, 0);
      write(32'h0003084C, 0);
      write(32'h00030850, 0);
      write(32'h00030854, 0);
      write(32'h00030858, 0);
      write(32'h0003085C, 0);
      write(32'h00030860, 163);
      write(32'h00030864, 255);
      write(32'h00030868, 124);
      write(32'h0003086C, 0);
      write(32'h00030870, 0);
      write(32'h00030874, 0);
      write(32'h00030878, 0);
      write(32'h0003087C, 0);
      write(32'h00030880, 51);
      write(32'h00030884, 37);
      write(32'h00030888, 0);
      write(32'h0003088C, 0);
      write(32'h00030890, 0);
      write(32'h00030894, 0);
      write(32'h00030898, 82);
      write(32'h0003089C, 255);
      write(32'h000308A0, 203);
      write(32'h000308A4, 9);
      write(32'h000308A8, 0);
      write(32'h000308AC, 0);
      write(32'h000308B0, 0);
      write(32'h000308B4, 0);
      write(32'h000308B8, 0);
      write(32'h000308BC, 0);
      write(32'h000308C0, 0);
      write(32'h000308C4, 0);
      write(32'h000308C8, 0);
      write(32'h000308CC, 0);
      write(32'h000308D0, 96);
      write(32'h000308D4, 255);
      write(32'h000308D8, 184);
      write(32'h000308DC, 4);
      write(32'h000308E0, 0);
      write(32'h000308E4, 0);
      write(32'h000308E8, 0);
      write(32'h000308EC, 0);
      write(32'h000308F0, 180);
      write(32'h000308F4, 233);
      write(32'h000308F8, 79);
      write(32'h000308FC, 0);
      write(32'h00030900, 0);
      write(32'h00030904, 0);
      write(32'h00030908, 56);
      write(32'h0003090C, 251);
      write(32'h00030910, 189);
      write(32'h00030914, 19);
      write(32'h00030918, 0);
      write(32'h0003091C, 0);
      write(32'h00030920, 0);
      write(32'h00030924, 0);
      write(32'h00030928, 0);
      write(32'h0003092C, 0);
      write(32'h00030930, 0);
      write(32'h00030934, 0);
      write(32'h00030938, 0);
      write(32'h0003093C, 0);
      write(32'h00030940, 31);
      write(32'h00030944, 235);
      write(32'h00030948, 236);
      write(32'h0003094C, 42);
      write(32'h00030950, 0);
      write(32'h00030954, 0);
      write(32'h00030958, 0);
      write(32'h0003095C, 42);
      write(32'h00030960, 238);
      write(32'h00030964, 252);
      write(32'h00030968, 64);
      write(32'h0003096C, 0);
      write(32'h00030970, 0);
      write(32'h00030974, 0);
      write(32'h00030978, 12);
      write(32'h0003097C, 61);
      write(32'h00030980, 29);
      write(32'h00030984, 2);
      write(32'h00030988, 0);
      write(32'h0003098C, 0);
      write(32'h00030990, 0);
      write(32'h00030994, 0);
      write(32'h00030998, 0);
      write(32'h0003099C, 0);
      write(32'h000309A0, 0);
      write(32'h000309A4, 0);
      write(32'h000309A8, 0);
      write(32'h000309AC, 0);
      write(32'h000309B0, 3);
      write(32'h000309B4, 162);
      write(32'h000309B8, 255);
      write(32'h000309BC, 121);
      write(32'h000309C0, 0);
      write(32'h000309C4, 0);
      write(32'h000309C8, 0);
      write(32'h000309CC, 133);
      write(32'h000309D0, 255);
      write(32'h000309D4, 168);
      write(32'h000309D8, 1);
      write(32'h000309DC, 0);
      write(32'h000309E0, 0);
      write(32'h000309E4, 0);
      write(32'h000309E8, 0);
      write(32'h000309EC, 0);
      write(32'h000309F0, 0);
      write(32'h000309F4, 0);
      write(32'h000309F8, 0);
      write(32'h000309FC, 0);
      write(32'h00030A00, 0);
      write(32'h00030A04, 0);
      write(32'h00030A08, 0);
      write(32'h00030A0C, 0);
      write(32'h00030A10, 0);
      write(32'h00030A14, 0);
      write(32'h00030A18, 0);
      write(32'h00030A1C, 0);
      write(32'h00030A20, 0);
      write(32'h00030A24, 65);
      write(32'h00030A28, 249);
      write(32'h00030A2C, 227);
      write(32'h00030A30, 29);
      write(32'h00030A34, 0);
      write(32'h00030A38, 39);
      write(32'h00030A3C, 235);
      write(32'h00030A40, 239);
      write(32'h00030A44, 50);
      write(32'h00030A48, 0);
      write(32'h00030A4C, 0);
      write(32'h00030A50, 0);
      write(32'h00030A54, 0);
      write(32'h00030A58, 0);
      write(32'h00030A5C, 0);
      write(32'h00030A60, 0);
      write(32'h00030A64, 0);
      write(32'h00030A68, 0);
      write(32'h00030A6C, 0);
      write(32'h00030A70, 0);
      write(32'h00030A74, 0);
      write(32'h00030A78, 0);
      write(32'h00030A7C, 0);
      write(32'h00030A80, 0);
      write(32'h00030A84, 0);
      write(32'h00030A88, 0);
      write(32'h00030A8C, 0);
      write(32'h00030A90, 0);
      write(32'h00030A94, 0);
      write(32'h00030A98, 161);
      write(32'h00030A9C, 255);
      write(32'h00030AA0, 174);
      write(32'h00030AA4, 53);
      write(32'h00030AA8, 185);
      write(32'h00030AAC, 255);
      write(32'h00030AB0, 125);
      write(32'h00030AB4, 0);
      write(32'h00030AB8, 0);
      write(32'h00030ABC, 0);
      write(32'h00030AC0, 0);
      write(32'h00030AC4, 0);
      write(32'h00030AC8, 0);
      write(32'h00030ACC, 0);
      write(32'h00030AD0, 0);
      write(32'h00030AD4, 0);
      write(32'h00030AD8, 0);
      write(32'h00030ADC, 0);
      write(32'h00030AE0, 0);
      write(32'h00030AE4, 0);
      write(32'h00030AE8, 0);
      write(32'h00030AEC, 0);
      write(32'h00030AF0, 0);
      write(32'h00030AF4, 0);
      write(32'h00030AF8, 0);
      write(32'h00030AFC, 0);
      write(32'h00030B00, 0);
      write(32'h00030B04, 0);
      write(32'h00030B08, 28);
      write(32'h00030B0C, 205);
      write(32'h00030B10, 255);
      write(32'h00030B14, 255);
      write(32'h00030B18, 255);
      write(32'h00030B1C, 165);
      write(32'h00030B20, 11);
      write(32'h00030B24, 0);
      write(32'h00030B28, 0);
      write(32'h00030B2C, 0);
      write(32'h00030B30, 0);
      write(32'h00030B34, 0);
      write(32'h00030B38, 0);
      write(32'h00030B3C, 0);
      write(32'h00030B40, 0);
      write(32'h00030B44, 0);
      write(32'h00030B48, 0);
      write(32'h00030B4C, 0);
      write(32'h00030B50, 0);
      write(32'h00030B54, 0);
      write(32'h00030B58, 0);
      write(32'h00030B5C, 0);
      write(32'h00030B60, 0);
      write(32'h00030B64, 0);
      write(32'h00030B68, 0);
      write(32'h00030B6C, 0);
      write(32'h00030B70, 0);
      write(32'h00030B74, 0);
      write(32'h00030B78, 0);
      write(32'h00030B7C, 30);
      write(32'h00030B80, 146);
      write(32'h00030B84, 192);
      write(32'h00030B88, 117);
      write(32'h00030B8C, 11);
      write(32'h00030B90, 0);
      write(32'h00030B94, 0);
      write(32'h00030B98, 0);
      write(32'h00030B9C, 0);
      write(32'h00030BA0, 0);
      write(32'h00030BA4, 0);
      write(32'h00030BA8, 0);
      write(32'h00030BAC, 0);
      write(32'h00030BB0, 0);
      write(32'h00030BB4, 0);
      write(32'h00030BB8, 0);
      write(32'h00030BBC, 0);
      write(32'h00030BC0, 0);
      write(32'h00030BC4, 0);
      write(32'h00030BC8, 0);
      write(32'h00030BCC, 0);
      write(32'h00030BD0, 0);
      write(32'h00030BD4, 0);
      write(32'h00030BD8, 0);
      write(32'h00030BDC, 0);
      write(32'h00030BE0, 0);
      write(32'h00030BE4, 0);
      write(32'h00030BE8, 0);
      write(32'h00030BEC, 0);
      write(32'h00030BF0, 0);
      write(32'h00030BF4, 0);
      write(32'h00030BF8, 0);
      write(32'h00030BFC, 0);
      write(32'h00030C00, 0);
      write(32'h00030C04, 0);
      write(32'h00030C08, 0);
      write(32'h00030C0C, 0);
      write(32'h00030C10, 0);
      write(32'h00030C14, 0);
      write(32'h00030C18, 0);
      write(32'h00030C1C, 0);
      write(32'h00030C20, 0);
      write(32'h00030C24, 0);
      write(32'h00030C28, 0);
      write(32'h00030C2C, 0);
      write(32'h00030C30, 0);
      write(32'h00030C34, 0);
      write(32'h00030C38, 0);
      write(32'h00030C3C, 0);


      $display("DATA I");


      
      #1000 $finish;
   end

   task write;
      input [31:0] adr_i;
      input [31:0] data_i;
      begin
	 WR = 1; ADR = adr_i; WDATA = data_i;
	 #(PERIOD)
	 WR = 0;
	 #(PERIOD);
      end
   endtask //
   
   
endmodule // sim_a_tb
