module img_sram
  (
   input 	    CLK,
   input 	    CS,
   input 	    WR,
   input [11:0]     ADR,
   input [7:0] 	    WDATA,
   output [28*28*8-1:0] RDATA
   
   );

   wire [9:0] 	    local_adr;

   assign local_adr = ADR[11:2];

   reg [7:0] 	    RDATA_00;
   reg [7:0] 	    RDATA_01;
   reg [7:0] 	    RDATA_02;
   reg [7:0] 	    RDATA_03;
   reg [7:0] 	    RDATA_04;
   reg [7:0] 	    RDATA_05;
   reg [7:0] 	    RDATA_06;
   reg [7:0] 	    RDATA_07;
   reg [7:0] 	    RDATA_08;
   reg [7:0] 	    RDATA_09;
   reg [7:0] 	    RDATA_10;
   reg [7:0] 	    RDATA_11;
   reg [7:0] 	    RDATA_12;
   reg [7:0] 	    RDATA_13;
   reg [7:0] 	    RDATA_14;
   reg [7:0] 	    RDATA_15;
   reg [7:0] 	    RDATA_16;
   reg [7:0] 	    RDATA_17;
   reg [7:0] 	    RDATA_18;
   reg [7:0] 	    RDATA_19;
   reg [7:0] 	    RDATA_20;
   reg [7:0] 	    RDATA_21;
   reg [7:0] 	    RDATA_22;
   reg [7:0] 	    RDATA_23;
   reg [7:0] 	    RDATA_24;
   reg [7:0] 	    RDATA_25;
   reg [7:0] 	    RDATA_26;
   reg [7:0] 	    RDATA_27;
   reg [7:0] 	    RDATA_28;
   reg [7:0] 	    RDATA_29;
   reg [7:0] 	    RDATA_30;
   reg [7:0] 	    RDATA_31;
   reg [7:0] 	    RDATA_32;
   reg [7:0] 	    RDATA_33;
   reg [7:0] 	    RDATA_34;
   reg [7:0] 	    RDATA_35;
   reg [7:0] 	    RDATA_36;
   reg [7:0] 	    RDATA_37;
   reg [7:0] 	    RDATA_38;
   reg [7:0] 	    RDATA_39;
   reg [7:0] 	    RDATA_40;
   reg [7:0] 	    RDATA_41;
   reg [7:0] 	    RDATA_42;
   reg [7:0] 	    RDATA_43;
   reg [7:0] 	    RDATA_44;
   reg [7:0] 	    RDATA_45;
   reg [7:0] 	    RDATA_46;
   reg [7:0] 	    RDATA_47;
   reg [7:0] 	    RDATA_48;
   reg [7:0] 	    RDATA_49;
   reg [7:0] 	    RDATA_50;
   reg [7:0] 	    RDATA_51;
   reg [7:0] 	    RDATA_52;
   reg [7:0] 	    RDATA_53;
   reg [7:0] 	    RDATA_54;
   reg [7:0] 	    RDATA_55;
   reg [7:0] 	    RDATA_56;
   reg [7:0] 	    RDATA_57;
   reg [7:0] 	    RDATA_58;
   reg [7:0] 	    RDATA_59;
   reg [7:0] 	    RDATA_60;
   reg [7:0] 	    RDATA_61;
   reg [7:0] 	    RDATA_62;
   reg [7:0] 	    RDATA_63;
   reg [7:0] 	    RDATA_64;
   reg [7:0] 	    RDATA_65;
   reg [7:0] 	    RDATA_66;
   reg [7:0] 	    RDATA_67;
   reg [7:0] 	    RDATA_68;
   reg [7:0] 	    RDATA_69;
   reg [7:0] 	    RDATA_70;
   reg [7:0] 	    RDATA_71;
   reg [7:0] 	    RDATA_72;
   reg [7:0] 	    RDATA_73;
   reg [7:0] 	    RDATA_74;
   reg [7:0] 	    RDATA_75;
   reg [7:0] 	    RDATA_76;
   reg [7:0] 	    RDATA_77;
   reg [7:0] 	    RDATA_78;
   reg [7:0] 	    RDATA_79;
   reg [7:0] 	    RDATA_80;
   reg [7:0] 	    RDATA_81;
   reg [7:0] 	    RDATA_82;
   reg [7:0] 	    RDATA_83;
   reg [7:0] 	    RDATA_84;
   reg [7:0] 	    RDATA_85;
   reg [7:0] 	    RDATA_86;
   reg [7:0] 	    RDATA_87;
   reg [7:0] 	    RDATA_88;
   reg [7:0] 	    RDATA_89;
   reg [7:0] 	    RDATA_90;
   reg [7:0] 	    RDATA_91;
   reg [7:0] 	    RDATA_92;
   reg [7:0] 	    RDATA_93;
   reg [7:0] 	    RDATA_94;
   reg [7:0] 	    RDATA_95;
   reg [7:0] 	    RDATA_96;
   reg [7:0] 	    RDATA_97;
   reg [7:0] 	    RDATA_98;
   reg [7:0] 	    RDATA_99;
   reg [7:0] 	    RDATA_100;
   reg [7:0] 	    RDATA_101;
   reg [7:0] 	    RDATA_102;
   reg [7:0] 	    RDATA_103;
   reg [7:0] 	    RDATA_104;
   reg [7:0] 	    RDATA_105;
   reg [7:0] 	    RDATA_106;
   reg [7:0] 	    RDATA_107;
   reg [7:0] 	    RDATA_108;
   reg [7:0] 	    RDATA_109;
   reg [7:0] 	    RDATA_110;
   reg [7:0] 	    RDATA_111;
   reg [7:0] 	    RDATA_112;
   reg [7:0] 	    RDATA_113;
   reg [7:0] 	    RDATA_114;
   reg [7:0] 	    RDATA_115;
   reg [7:0] 	    RDATA_116;
   reg [7:0] 	    RDATA_117;
   reg [7:0] 	    RDATA_118;
   reg [7:0] 	    RDATA_119;
   reg [7:0] 	    RDATA_120;
   reg [7:0] 	    RDATA_121;
   reg [7:0] 	    RDATA_122;
   reg [7:0] 	    RDATA_123;
   reg [7:0] 	    RDATA_124;
   reg [7:0] 	    RDATA_125;
   reg [7:0] 	    RDATA_126;
   reg [7:0] 	    RDATA_127;
   reg [7:0] 	    RDATA_128;
   reg [7:0] 	    RDATA_129;
   reg [7:0] 	    RDATA_130;
   reg [7:0] 	    RDATA_131;
   reg [7:0] 	    RDATA_132;
   reg [7:0] 	    RDATA_133;
   reg [7:0] 	    RDATA_134;
   reg [7:0] 	    RDATA_135;
   reg [7:0] 	    RDATA_136;
   reg [7:0] 	    RDATA_137;
   reg [7:0] 	    RDATA_138;
   reg [7:0] 	    RDATA_139;
   reg [7:0] 	    RDATA_140;
   reg [7:0] 	    RDATA_141;
   reg [7:0] 	    RDATA_142;
   reg [7:0] 	    RDATA_143;
   reg [7:0] 	    RDATA_144;
   reg [7:0] 	    RDATA_145;
   reg [7:0] 	    RDATA_146;
   reg [7:0] 	    RDATA_147;
   reg [7:0] 	    RDATA_148;
   reg [7:0] 	    RDATA_149;
   reg [7:0] 	    RDATA_150;
   reg [7:0] 	    RDATA_151;
   reg [7:0] 	    RDATA_152;
   reg [7:0] 	    RDATA_153;
   reg [7:0] 	    RDATA_154;
   reg [7:0] 	    RDATA_155;
   reg [7:0] 	    RDATA_156;
   reg [7:0] 	    RDATA_157;
   reg [7:0] 	    RDATA_158;
   reg [7:0] 	    RDATA_159;
   reg [7:0] 	    RDATA_160;
   reg [7:0] 	    RDATA_161;
   reg [7:0] 	    RDATA_162;
   reg [7:0] 	    RDATA_163;
   reg [7:0] 	    RDATA_164;
   reg [7:0] 	    RDATA_165;
   reg [7:0] 	    RDATA_166;
   reg [7:0] 	    RDATA_167;
   reg [7:0] 	    RDATA_168;
   reg [7:0] 	    RDATA_169;
   reg [7:0] 	    RDATA_170;
   reg [7:0] 	    RDATA_171;
   reg [7:0] 	    RDATA_172;
   reg [7:0] 	    RDATA_173;
   reg [7:0] 	    RDATA_174;
   reg [7:0] 	    RDATA_175;
   reg [7:0] 	    RDATA_176;
   reg [7:0] 	    RDATA_177;
   reg [7:0] 	    RDATA_178;
   reg [7:0] 	    RDATA_179;
   reg [7:0] 	    RDATA_180;
   reg [7:0] 	    RDATA_181;
   reg [7:0] 	    RDATA_182;
   reg [7:0] 	    RDATA_183;
   reg [7:0] 	    RDATA_184;
   reg [7:0] 	    RDATA_185;
   reg [7:0] 	    RDATA_186;
   reg [7:0] 	    RDATA_187;
   reg [7:0] 	    RDATA_188;
   reg [7:0] 	    RDATA_189;
   reg [7:0] 	    RDATA_190;
   reg [7:0] 	    RDATA_191;
   reg [7:0] 	    RDATA_192;
   reg [7:0] 	    RDATA_193;
   reg [7:0] 	    RDATA_194;
   reg [7:0] 	    RDATA_195;
   reg [7:0] 	    RDATA_196;
   reg [7:0] 	    RDATA_197;
   reg [7:0] 	    RDATA_198;
   reg [7:0] 	    RDATA_199;
   reg [7:0] 	    RDATA_200;
   reg [7:0] 	    RDATA_201;
   reg [7:0] 	    RDATA_202;
   reg [7:0] 	    RDATA_203;
   reg [7:0] 	    RDATA_204;
   reg [7:0] 	    RDATA_205;
   reg [7:0] 	    RDATA_206;
   reg [7:0] 	    RDATA_207;
   reg [7:0] 	    RDATA_208;
   reg [7:0] 	    RDATA_209;
   reg [7:0] 	    RDATA_210;
   reg [7:0] 	    RDATA_211;
   reg [7:0] 	    RDATA_212;
   reg [7:0] 	    RDATA_213;
   reg [7:0] 	    RDATA_214;
   reg [7:0] 	    RDATA_215;
   reg [7:0] 	    RDATA_216;
   reg [7:0] 	    RDATA_217;
   reg [7:0] 	    RDATA_218;
   reg [7:0] 	    RDATA_219;
   reg [7:0] 	    RDATA_220;
   reg [7:0] 	    RDATA_221;
   reg [7:0] 	    RDATA_222;
   reg [7:0] 	    RDATA_223;
   reg [7:0] 	    RDATA_224;
   reg [7:0] 	    RDATA_225;
   reg [7:0] 	    RDATA_226;
   reg [7:0] 	    RDATA_227;
   reg [7:0] 	    RDATA_228;
   reg [7:0] 	    RDATA_229;
   reg [7:0] 	    RDATA_230;
   reg [7:0] 	    RDATA_231;
   reg [7:0] 	    RDATA_232;
   reg [7:0] 	    RDATA_233;
   reg [7:0] 	    RDATA_234;
   reg [7:0] 	    RDATA_235;
   reg [7:0] 	    RDATA_236;
   reg [7:0] 	    RDATA_237;
   reg [7:0] 	    RDATA_238;
   reg [7:0] 	    RDATA_239;
   reg [7:0] 	    RDATA_240;
   reg [7:0] 	    RDATA_241;
   reg [7:0] 	    RDATA_242;
   reg [7:0] 	    RDATA_243;
   reg [7:0] 	    RDATA_244;
   reg [7:0] 	    RDATA_245;
   reg [7:0] 	    RDATA_246;
   reg [7:0] 	    RDATA_247;
   reg [7:0] 	    RDATA_248;
   reg [7:0] 	    RDATA_249;
   reg [7:0] 	    RDATA_250;
   reg [7:0] 	    RDATA_251;
   reg [7:0] 	    RDATA_252;
   reg [7:0] 	    RDATA_253;
   reg [7:0] 	    RDATA_254;
   reg [7:0] 	    RDATA_255;
   reg [7:0] 	    RDATA_256;
   reg [7:0] 	    RDATA_257;
   reg [7:0] 	    RDATA_258;
   reg [7:0] 	    RDATA_259;
   reg [7:0] 	    RDATA_260;
   reg [7:0] 	    RDATA_261;
   reg [7:0] 	    RDATA_262;
   reg [7:0] 	    RDATA_263;
   reg [7:0] 	    RDATA_264;
   reg [7:0] 	    RDATA_265;
   reg [7:0] 	    RDATA_266;
   reg [7:0] 	    RDATA_267;
   reg [7:0] 	    RDATA_268;
   reg [7:0] 	    RDATA_269;
   reg [7:0] 	    RDATA_270;
   reg [7:0] 	    RDATA_271;
   reg [7:0] 	    RDATA_272;
   reg [7:0] 	    RDATA_273;
   reg [7:0] 	    RDATA_274;
   reg [7:0] 	    RDATA_275;
   reg [7:0] 	    RDATA_276;
   reg [7:0] 	    RDATA_277;
   reg [7:0] 	    RDATA_278;
   reg [7:0] 	    RDATA_279;
   reg [7:0] 	    RDATA_280;
   reg [7:0] 	    RDATA_281;
   reg [7:0] 	    RDATA_282;
   reg [7:0] 	    RDATA_283;
   reg [7:0] 	    RDATA_284;
   reg [7:0] 	    RDATA_285;
   reg [7:0] 	    RDATA_286;
   reg [7:0] 	    RDATA_287;
   reg [7:0] 	    RDATA_288;
   reg [7:0] 	    RDATA_289;
   reg [7:0] 	    RDATA_290;
   reg [7:0] 	    RDATA_291;
   reg [7:0] 	    RDATA_292;
   reg [7:0] 	    RDATA_293;
   reg [7:0] 	    RDATA_294;
   reg [7:0] 	    RDATA_295;
   reg [7:0] 	    RDATA_296;
   reg [7:0] 	    RDATA_297;
   reg [7:0] 	    RDATA_298;
   reg [7:0] 	    RDATA_299;
   reg [7:0] 	    RDATA_300;
   reg [7:0] 	    RDATA_301;
   reg [7:0] 	    RDATA_302;
   reg [7:0] 	    RDATA_303;
   reg [7:0] 	    RDATA_304;
   reg [7:0] 	    RDATA_305;
   reg [7:0] 	    RDATA_306;
   reg [7:0] 	    RDATA_307;
   reg [7:0] 	    RDATA_308;
   reg [7:0] 	    RDATA_309;
   reg [7:0] 	    RDATA_310;
   reg [7:0] 	    RDATA_311;
   reg [7:0] 	    RDATA_312;
   reg [7:0] 	    RDATA_313;
   reg [7:0] 	    RDATA_314;
   reg [7:0] 	    RDATA_315;
   reg [7:0] 	    RDATA_316;
   reg [7:0] 	    RDATA_317;
   reg [7:0] 	    RDATA_318;
   reg [7:0] 	    RDATA_319;
   reg [7:0] 	    RDATA_320;
   reg [7:0] 	    RDATA_321;
   reg [7:0] 	    RDATA_322;
   reg [7:0] 	    RDATA_323;
   reg [7:0] 	    RDATA_324;
   reg [7:0] 	    RDATA_325;
   reg [7:0] 	    RDATA_326;
   reg [7:0] 	    RDATA_327;
   reg [7:0] 	    RDATA_328;
   reg [7:0] 	    RDATA_329;
   reg [7:0] 	    RDATA_330;
   reg [7:0] 	    RDATA_331;
   reg [7:0] 	    RDATA_332;
   reg [7:0] 	    RDATA_333;
   reg [7:0] 	    RDATA_334;
   reg [7:0] 	    RDATA_335;
   reg [7:0] 	    RDATA_336;
   reg [7:0] 	    RDATA_337;
   reg [7:0] 	    RDATA_338;
   reg [7:0] 	    RDATA_339;
   reg [7:0] 	    RDATA_340;
   reg [7:0] 	    RDATA_341;
   reg [7:0] 	    RDATA_342;
   reg [7:0] 	    RDATA_343;
   reg [7:0] 	    RDATA_344;
   reg [7:0] 	    RDATA_345;
   reg [7:0] 	    RDATA_346;
   reg [7:0] 	    RDATA_347;
   reg [7:0] 	    RDATA_348;
   reg [7:0] 	    RDATA_349;
   reg [7:0] 	    RDATA_350;
   reg [7:0] 	    RDATA_351;
   reg [7:0] 	    RDATA_352;
   reg [7:0] 	    RDATA_353;
   reg [7:0] 	    RDATA_354;
   reg [7:0] 	    RDATA_355;
   reg [7:0] 	    RDATA_356;
   reg [7:0] 	    RDATA_357;
   reg [7:0] 	    RDATA_358;
   reg [7:0] 	    RDATA_359;
   reg [7:0] 	    RDATA_360;
   reg [7:0] 	    RDATA_361;
   reg [7:0] 	    RDATA_362;
   reg [7:0] 	    RDATA_363;
   reg [7:0] 	    RDATA_364;
   reg [7:0] 	    RDATA_365;
   reg [7:0] 	    RDATA_366;
   reg [7:0] 	    RDATA_367;
   reg [7:0] 	    RDATA_368;
   reg [7:0] 	    RDATA_369;
   reg [7:0] 	    RDATA_370;
   reg [7:0] 	    RDATA_371;
   reg [7:0] 	    RDATA_372;
   reg [7:0] 	    RDATA_373;
   reg [7:0] 	    RDATA_374;
   reg [7:0] 	    RDATA_375;
   reg [7:0] 	    RDATA_376;
   reg [7:0] 	    RDATA_377;
   reg [7:0] 	    RDATA_378;
   reg [7:0] 	    RDATA_379;
   reg [7:0] 	    RDATA_380;
   reg [7:0] 	    RDATA_381;
   reg [7:0] 	    RDATA_382;
   reg [7:0] 	    RDATA_383;
   reg [7:0] 	    RDATA_384;
   reg [7:0] 	    RDATA_385;
   reg [7:0] 	    RDATA_386;
   reg [7:0] 	    RDATA_387;
   reg [7:0] 	    RDATA_388;
   reg [7:0] 	    RDATA_389;
   reg [7:0] 	    RDATA_390;
   reg [7:0] 	    RDATA_391;
   reg [7:0] 	    RDATA_392;
   reg [7:0] 	    RDATA_393;
   reg [7:0] 	    RDATA_394;
   reg [7:0] 	    RDATA_395;
   reg [7:0] 	    RDATA_396;
   reg [7:0] 	    RDATA_397;
   reg [7:0] 	    RDATA_398;
   reg [7:0] 	    RDATA_399;
   reg [7:0] 	    RDATA_400;
   reg [7:0] 	    RDATA_401;
   reg [7:0] 	    RDATA_402;
   reg [7:0] 	    RDATA_403;
   reg [7:0] 	    RDATA_404;
   reg [7:0] 	    RDATA_405;
   reg [7:0] 	    RDATA_406;
   reg [7:0] 	    RDATA_407;
   reg [7:0] 	    RDATA_408;
   reg [7:0] 	    RDATA_409;
   reg [7:0] 	    RDATA_410;
   reg [7:0] 	    RDATA_411;
   reg [7:0] 	    RDATA_412;
   reg [7:0] 	    RDATA_413;
   reg [7:0] 	    RDATA_414;
   reg [7:0] 	    RDATA_415;
   reg [7:0] 	    RDATA_416;
   reg [7:0] 	    RDATA_417;
   reg [7:0] 	    RDATA_418;
   reg [7:0] 	    RDATA_419;
   reg [7:0] 	    RDATA_420;
   reg [7:0] 	    RDATA_421;
   reg [7:0] 	    RDATA_422;
   reg [7:0] 	    RDATA_423;
   reg [7:0] 	    RDATA_424;
   reg [7:0] 	    RDATA_425;
   reg [7:0] 	    RDATA_426;
   reg [7:0] 	    RDATA_427;
   reg [7:0] 	    RDATA_428;
   reg [7:0] 	    RDATA_429;
   reg [7:0] 	    RDATA_430;
   reg [7:0] 	    RDATA_431;
   reg [7:0] 	    RDATA_432;
   reg [7:0] 	    RDATA_433;
   reg [7:0] 	    RDATA_434;
   reg [7:0] 	    RDATA_435;
   reg [7:0] 	    RDATA_436;
   reg [7:0] 	    RDATA_437;
   reg [7:0] 	    RDATA_438;
   reg [7:0] 	    RDATA_439;
   reg [7:0] 	    RDATA_440;
   reg [7:0] 	    RDATA_441;
   reg [7:0] 	    RDATA_442;
   reg [7:0] 	    RDATA_443;
   reg [7:0] 	    RDATA_444;
   reg [7:0] 	    RDATA_445;
   reg [7:0] 	    RDATA_446;
   reg [7:0] 	    RDATA_447;
   reg [7:0] 	    RDATA_448;
   reg [7:0] 	    RDATA_449;
   reg [7:0] 	    RDATA_450;
   reg [7:0] 	    RDATA_451;
   reg [7:0] 	    RDATA_452;
   reg [7:0] 	    RDATA_453;
   reg [7:0] 	    RDATA_454;
   reg [7:0] 	    RDATA_455;
   reg [7:0] 	    RDATA_456;
   reg [7:0] 	    RDATA_457;
   reg [7:0] 	    RDATA_458;
   reg [7:0] 	    RDATA_459;
   reg [7:0] 	    RDATA_460;
   reg [7:0] 	    RDATA_461;
   reg [7:0] 	    RDATA_462;
   reg [7:0] 	    RDATA_463;
   reg [7:0] 	    RDATA_464;
   reg [7:0] 	    RDATA_465;
   reg [7:0] 	    RDATA_466;
   reg [7:0] 	    RDATA_467;
   reg [7:0] 	    RDATA_468;
   reg [7:0] 	    RDATA_469;
   reg [7:0] 	    RDATA_470;
   reg [7:0] 	    RDATA_471;
   reg [7:0] 	    RDATA_472;
   reg [7:0] 	    RDATA_473;
   reg [7:0] 	    RDATA_474;
   reg [7:0] 	    RDATA_475;
   reg [7:0] 	    RDATA_476;
   reg [7:0] 	    RDATA_477;
   reg [7:0] 	    RDATA_478;
   reg [7:0] 	    RDATA_479;
   reg [7:0] 	    RDATA_480;
   reg [7:0] 	    RDATA_481;
   reg [7:0] 	    RDATA_482;
   reg [7:0] 	    RDATA_483;
   reg [7:0] 	    RDATA_484;
   reg [7:0] 	    RDATA_485;
   reg [7:0] 	    RDATA_486;
   reg [7:0] 	    RDATA_487;
   reg [7:0] 	    RDATA_488;
   reg [7:0] 	    RDATA_489;
   reg [7:0] 	    RDATA_490;
   reg [7:0] 	    RDATA_491;
   reg [7:0] 	    RDATA_492;
   reg [7:0] 	    RDATA_493;
   reg [7:0] 	    RDATA_494;
   reg [7:0] 	    RDATA_495;
   reg [7:0] 	    RDATA_496;
   reg [7:0] 	    RDATA_497;
   reg [7:0] 	    RDATA_498;
   reg [7:0] 	    RDATA_499;
   reg [7:0] 	    RDATA_500;
   reg [7:0] 	    RDATA_501;
   reg [7:0] 	    RDATA_502;
   reg [7:0] 	    RDATA_503;
   reg [7:0] 	    RDATA_504;
   reg [7:0] 	    RDATA_505;
   reg [7:0] 	    RDATA_506;
   reg [7:0] 	    RDATA_507;
   reg [7:0] 	    RDATA_508;
   reg [7:0] 	    RDATA_509;
   reg [7:0] 	    RDATA_510;
   reg [7:0] 	    RDATA_511;
   reg [7:0] 	    RDATA_512;
   reg [7:0] 	    RDATA_513;
   reg [7:0] 	    RDATA_514;
   reg [7:0] 	    RDATA_515;
   reg [7:0] 	    RDATA_516;
   reg [7:0] 	    RDATA_517;
   reg [7:0] 	    RDATA_518;
   reg [7:0] 	    RDATA_519;
   reg [7:0] 	    RDATA_520;
   reg [7:0] 	    RDATA_521;
   reg [7:0] 	    RDATA_522;
   reg [7:0] 	    RDATA_523;
   reg [7:0] 	    RDATA_524;
   reg [7:0] 	    RDATA_525;
   reg [7:0] 	    RDATA_526;
   reg [7:0] 	    RDATA_527;
   reg [7:0] 	    RDATA_528;
   reg [7:0] 	    RDATA_529;
   reg [7:0] 	    RDATA_530;
   reg [7:0] 	    RDATA_531;
   reg [7:0] 	    RDATA_532;
   reg [7:0] 	    RDATA_533;
   reg [7:0] 	    RDATA_534;
   reg [7:0] 	    RDATA_535;
   reg [7:0] 	    RDATA_536;
   reg [7:0] 	    RDATA_537;
   reg [7:0] 	    RDATA_538;
   reg [7:0] 	    RDATA_539;
   reg [7:0] 	    RDATA_540;
   reg [7:0] 	    RDATA_541;
   reg [7:0] 	    RDATA_542;
   reg [7:0] 	    RDATA_543;
   reg [7:0] 	    RDATA_544;
   reg [7:0] 	    RDATA_545;
   reg [7:0] 	    RDATA_546;
   reg [7:0] 	    RDATA_547;
   reg [7:0] 	    RDATA_548;
   reg [7:0] 	    RDATA_549;
   reg [7:0] 	    RDATA_550;
   reg [7:0] 	    RDATA_551;
   reg [7:0] 	    RDATA_552;
   reg [7:0] 	    RDATA_553;
   reg [7:0] 	    RDATA_554;
   reg [7:0] 	    RDATA_555;
   reg [7:0] 	    RDATA_556;
   reg [7:0] 	    RDATA_557;
   reg [7:0] 	    RDATA_558;
   reg [7:0] 	    RDATA_559;
   reg [7:0] 	    RDATA_560;
   reg [7:0] 	    RDATA_561;
   reg [7:0] 	    RDATA_562;
   reg [7:0] 	    RDATA_563;
   reg [7:0] 	    RDATA_564;
   reg [7:0] 	    RDATA_565;
   reg [7:0] 	    RDATA_566;
   reg [7:0] 	    RDATA_567;
   reg [7:0] 	    RDATA_568;
   reg [7:0] 	    RDATA_569;
   reg [7:0] 	    RDATA_570;
   reg [7:0] 	    RDATA_571;
   reg [7:0] 	    RDATA_572;
   reg [7:0] 	    RDATA_573;
   reg [7:0] 	    RDATA_574;
   reg [7:0] 	    RDATA_575;
   reg [7:0] 	    RDATA_576;
   reg [7:0] 	    RDATA_577;
   reg [7:0] 	    RDATA_578;
   reg [7:0] 	    RDATA_579;
   reg [7:0] 	    RDATA_580;
   reg [7:0] 	    RDATA_581;
   reg [7:0] 	    RDATA_582;
   reg [7:0] 	    RDATA_583;
   reg [7:0] 	    RDATA_584;
   reg [7:0] 	    RDATA_585;
   reg [7:0] 	    RDATA_586;
   reg [7:0] 	    RDATA_587;
   reg [7:0] 	    RDATA_588;
   reg [7:0] 	    RDATA_589;
   reg [7:0] 	    RDATA_590;
   reg [7:0] 	    RDATA_591;
   reg [7:0] 	    RDATA_592;
   reg [7:0] 	    RDATA_593;
   reg [7:0] 	    RDATA_594;
   reg [7:0] 	    RDATA_595;
   reg [7:0] 	    RDATA_596;
   reg [7:0] 	    RDATA_597;
   reg [7:0] 	    RDATA_598;
   reg [7:0] 	    RDATA_599;
   reg [7:0] 	    RDATA_600;
   reg [7:0] 	    RDATA_601;
   reg [7:0] 	    RDATA_602;
   reg [7:0] 	    RDATA_603;
   reg [7:0] 	    RDATA_604;
   reg [7:0] 	    RDATA_605;
   reg [7:0] 	    RDATA_606;
   reg [7:0] 	    RDATA_607;
   reg [7:0] 	    RDATA_608;
   reg [7:0] 	    RDATA_609;
   reg [7:0] 	    RDATA_610;
   reg [7:0] 	    RDATA_611;
   reg [7:0] 	    RDATA_612;
   reg [7:0] 	    RDATA_613;
   reg [7:0] 	    RDATA_614;
   reg [7:0] 	    RDATA_615;
   reg [7:0] 	    RDATA_616;
   reg [7:0] 	    RDATA_617;
   reg [7:0] 	    RDATA_618;
   reg [7:0] 	    RDATA_619;
   reg [7:0] 	    RDATA_620;
   reg [7:0] 	    RDATA_621;
   reg [7:0] 	    RDATA_622;
   reg [7:0] 	    RDATA_623;
   reg [7:0] 	    RDATA_624;
   reg [7:0] 	    RDATA_625;
   reg [7:0] 	    RDATA_626;
   reg [7:0] 	    RDATA_627;
   reg [7:0] 	    RDATA_628;
   reg [7:0] 	    RDATA_629;
   reg [7:0] 	    RDATA_630;
   reg [7:0] 	    RDATA_631;
   reg [7:0] 	    RDATA_632;
   reg [7:0] 	    RDATA_633;
   reg [7:0] 	    RDATA_634;
   reg [7:0] 	    RDATA_635;
   reg [7:0] 	    RDATA_636;
   reg [7:0] 	    RDATA_637;
   reg [7:0] 	    RDATA_638;
   reg [7:0] 	    RDATA_639;
   reg [7:0] 	    RDATA_640;
   reg [7:0] 	    RDATA_641;
   reg [7:0] 	    RDATA_642;
   reg [7:0] 	    RDATA_643;
   reg [7:0] 	    RDATA_644;
   reg [7:0] 	    RDATA_645;
   reg [7:0] 	    RDATA_646;
   reg [7:0] 	    RDATA_647;
   reg [7:0] 	    RDATA_648;
   reg [7:0] 	    RDATA_649;
   reg [7:0] 	    RDATA_650;
   reg [7:0] 	    RDATA_651;
   reg [7:0] 	    RDATA_652;
   reg [7:0] 	    RDATA_653;
   reg [7:0] 	    RDATA_654;
   reg [7:0] 	    RDATA_655;
   reg [7:0] 	    RDATA_656;
   reg [7:0] 	    RDATA_657;
   reg [7:0] 	    RDATA_658;
   reg [7:0] 	    RDATA_659;
   reg [7:0] 	    RDATA_660;
   reg [7:0] 	    RDATA_661;
   reg [7:0] 	    RDATA_662;
   reg [7:0] 	    RDATA_663;
   reg [7:0] 	    RDATA_664;
   reg [7:0] 	    RDATA_665;
   reg [7:0] 	    RDATA_666;
   reg [7:0] 	    RDATA_667;
   reg [7:0] 	    RDATA_668;
   reg [7:0] 	    RDATA_669;
   reg [7:0] 	    RDATA_670;
   reg [7:0] 	    RDATA_671;
   reg [7:0] 	    RDATA_672;
   reg [7:0] 	    RDATA_673;
   reg [7:0] 	    RDATA_674;
   reg [7:0] 	    RDATA_675;
   reg [7:0] 	    RDATA_676;
   reg [7:0] 	    RDATA_677;
   reg [7:0] 	    RDATA_678;
   reg [7:0] 	    RDATA_679;
   reg [7:0] 	    RDATA_680;
   reg [7:0] 	    RDATA_681;
   reg [7:0] 	    RDATA_682;
   reg [7:0] 	    RDATA_683;
   reg [7:0] 	    RDATA_684;
   reg [7:0] 	    RDATA_685;
   reg [7:0] 	    RDATA_686;
   reg [7:0] 	    RDATA_687;
   reg [7:0] 	    RDATA_688;
   reg [7:0] 	    RDATA_689;
   reg [7:0] 	    RDATA_690;
   reg [7:0] 	    RDATA_691;
   reg [7:0] 	    RDATA_692;
   reg [7:0] 	    RDATA_693;
   reg [7:0] 	    RDATA_694;
   reg [7:0] 	    RDATA_695;
   reg [7:0] 	    RDATA_696;
   reg [7:0] 	    RDATA_697;
   reg [7:0] 	    RDATA_698;
   reg [7:0] 	    RDATA_699;
   reg [7:0] 	    RDATA_700;
   reg [7:0] 	    RDATA_701;
   reg [7:0] 	    RDATA_702;
   reg [7:0] 	    RDATA_703;
   reg [7:0] 	    RDATA_704;
   reg [7:0] 	    RDATA_705;
   reg [7:0] 	    RDATA_706;
   reg [7:0] 	    RDATA_707;
   reg [7:0] 	    RDATA_708;
   reg [7:0] 	    RDATA_709;
   reg [7:0] 	    RDATA_710;
   reg [7:0] 	    RDATA_711;
   reg [7:0] 	    RDATA_712;
   reg [7:0] 	    RDATA_713;
   reg [7:0] 	    RDATA_714;
   reg [7:0] 	    RDATA_715;
   reg [7:0] 	    RDATA_716;
   reg [7:0] 	    RDATA_717;
   reg [7:0] 	    RDATA_718;
   reg [7:0] 	    RDATA_719;
   reg [7:0] 	    RDATA_720;
   reg [7:0] 	    RDATA_721;
   reg [7:0] 	    RDATA_722;
   reg [7:0] 	    RDATA_723;
   reg [7:0] 	    RDATA_724;
   reg [7:0] 	    RDATA_725;
   reg [7:0] 	    RDATA_726;
   reg [7:0] 	    RDATA_727;
   reg [7:0] 	    RDATA_728;
   reg [7:0] 	    RDATA_729;
   reg [7:0] 	    RDATA_730;
   reg [7:0] 	    RDATA_731;
   reg [7:0] 	    RDATA_732;
   reg [7:0] 	    RDATA_733;
   reg [7:0] 	    RDATA_734;
   reg [7:0] 	    RDATA_735;
   reg [7:0] 	    RDATA_736;
   reg [7:0] 	    RDATA_737;
   reg [7:0] 	    RDATA_738;
   reg [7:0] 	    RDATA_739;
   reg [7:0] 	    RDATA_740;
   reg [7:0] 	    RDATA_741;
   reg [7:0] 	    RDATA_742;
   reg [7:0] 	    RDATA_743;
   reg [7:0] 	    RDATA_744;
   reg [7:0] 	    RDATA_745;
   reg [7:0] 	    RDATA_746;
   reg [7:0] 	    RDATA_747;
   reg [7:0] 	    RDATA_748;
   reg [7:0] 	    RDATA_749;
   reg [7:0] 	    RDATA_750;
   reg [7:0] 	    RDATA_751;
   reg [7:0] 	    RDATA_752;
   reg [7:0] 	    RDATA_753;
   reg [7:0] 	    RDATA_754;
   reg [7:0] 	    RDATA_755;
   reg [7:0] 	    RDATA_756;
   reg [7:0] 	    RDATA_757;
   reg [7:0] 	    RDATA_758;
   reg [7:0] 	    RDATA_759;
   reg [7:0] 	    RDATA_760;
   reg [7:0] 	    RDATA_761;
   reg [7:0] 	    RDATA_762;
   reg [7:0] 	    RDATA_763;
   reg [7:0] 	    RDATA_764;
   reg [7:0] 	    RDATA_765;
   reg [7:0] 	    RDATA_766;
   reg [7:0] 	    RDATA_767;
   reg [7:0] 	    RDATA_768;
   reg [7:0] 	    RDATA_769;
   reg [7:0] 	    RDATA_770;
   reg [7:0] 	    RDATA_771;
   reg [7:0] 	    RDATA_772;
   reg [7:0] 	    RDATA_773;
   reg [7:0] 	    RDATA_774;
   reg [7:0] 	    RDATA_775;
   reg [7:0] 	    RDATA_776;
   reg [7:0] 	    RDATA_777;
   reg [7:0] 	    RDATA_778;
   reg [7:0] 	    RDATA_779;
   reg [7:0] 	    RDATA_780;
   reg [7:0] 	    RDATA_781;
   reg [7:0] 	    RDATA_782;
   reg [7:0] 	    RDATA_783;
   

   always @ (posedge CLK) begin
      if((CS == 1) & (WR == 1)) begin
	 if(local_adr==0) RDATA_00 <= WDATA;
	 if(local_adr==1) RDATA_01 <= WDATA;
	 if(local_adr==2) RDATA_02 <= WDATA;
	 if(local_adr==3) RDATA_03 <= WDATA;
	 if(local_adr==4) RDATA_04 <= WDATA;
	 if(local_adr==5) RDATA_05 <= WDATA;
	 if(local_adr==6) RDATA_06 <= WDATA;
	 if(local_adr==7) RDATA_07 <= WDATA;
	 if(local_adr==8) RDATA_08 <= WDATA;
	 if(local_adr==9) RDATA_09 <= WDATA;
	 if(local_adr==10) RDATA_10 <= WDATA;
	 if(local_adr==11) RDATA_11 <= WDATA;
	 if(local_adr==12) RDATA_12 <= WDATA;
	 if(local_adr==13) RDATA_13 <= WDATA;
	 if(local_adr==14) RDATA_14 <= WDATA;
	 if(local_adr==15) RDATA_15 <= WDATA;
	 if(local_adr==16) RDATA_16 <= WDATA;
	 if(local_adr==17) RDATA_17 <= WDATA;
	 if(local_adr==18) RDATA_18 <= WDATA;
	 if(local_adr==19) RDATA_19 <= WDATA;
	 if(local_adr==20) RDATA_20 <= WDATA;
	 if(local_adr==21) RDATA_21 <= WDATA;
	 if(local_adr==22) RDATA_22 <= WDATA;
	 if(local_adr==23) RDATA_23 <= WDATA;
	 if(local_adr==24) RDATA_24 <= WDATA;
	 if(local_adr==25) RDATA_25 <= WDATA;
	 if(local_adr==26) RDATA_26 <= WDATA;
	 if(local_adr==27) RDATA_27 <= WDATA;
	 if(local_adr==28) RDATA_28 <= WDATA;
	 if(local_adr==29) RDATA_29 <= WDATA;
	 if(local_adr==30) RDATA_30 <= WDATA;
	 if(local_adr==31) RDATA_31 <= WDATA;
	 if(local_adr==32) RDATA_32 <= WDATA;
	 if(local_adr==33) RDATA_33 <= WDATA;
	 if(local_adr==34) RDATA_34 <= WDATA;
	 if(local_adr==35) RDATA_35 <= WDATA;
	 if(local_adr==36) RDATA_36 <= WDATA;
	 if(local_adr==37) RDATA_37 <= WDATA;
	 if(local_adr==38) RDATA_38 <= WDATA;
	 if(local_adr==39) RDATA_39 <= WDATA;
	 if(local_adr==40) RDATA_40 <= WDATA;
	 if(local_adr==41) RDATA_41 <= WDATA;
	 if(local_adr==42) RDATA_42 <= WDATA;
	 if(local_adr==43) RDATA_43 <= WDATA;
	 if(local_adr==44) RDATA_44 <= WDATA;
	 if(local_adr==45) RDATA_45 <= WDATA;
	 if(local_adr==46) RDATA_46 <= WDATA;
	 if(local_adr==47) RDATA_47 <= WDATA;
	 if(local_adr==48) RDATA_48 <= WDATA;
	 if(local_adr==49) RDATA_49 <= WDATA;
	 if(local_adr==50) RDATA_50 <= WDATA;
	 if(local_adr==51) RDATA_51 <= WDATA;
	 if(local_adr==52) RDATA_52 <= WDATA;
	 if(local_adr==53) RDATA_53 <= WDATA;
	 if(local_adr==54) RDATA_54 <= WDATA;
	 if(local_adr==55) RDATA_55 <= WDATA;
	 if(local_adr==56) RDATA_56 <= WDATA;
	 if(local_adr==57) RDATA_57 <= WDATA;
	 if(local_adr==58) RDATA_58 <= WDATA;
	 if(local_adr==59) RDATA_59 <= WDATA;
	 if(local_adr==60) RDATA_60 <= WDATA;
	 if(local_adr==61) RDATA_61 <= WDATA;
	 if(local_adr==62) RDATA_62 <= WDATA;
	 if(local_adr==63) RDATA_63 <= WDATA;
	 if(local_adr==64) RDATA_64 <= WDATA;
	 if(local_adr==65) RDATA_65 <= WDATA;
	 if(local_adr==66) RDATA_66 <= WDATA;
	 if(local_adr==67) RDATA_67 <= WDATA;
	 if(local_adr==68) RDATA_68 <= WDATA;
	 if(local_adr==69) RDATA_69 <= WDATA;
	 if(local_adr==70) RDATA_70 <= WDATA;
	 if(local_adr==71) RDATA_71 <= WDATA;
	 if(local_adr==72) RDATA_72 <= WDATA;
	 if(local_adr==73) RDATA_73 <= WDATA;
	 if(local_adr==74) RDATA_74 <= WDATA;
	 if(local_adr==75) RDATA_75 <= WDATA;
	 if(local_adr==76) RDATA_76 <= WDATA;
	 if(local_adr==77) RDATA_77 <= WDATA;
	 if(local_adr==78) RDATA_78 <= WDATA;
	 if(local_adr==79) RDATA_79 <= WDATA;
	 if(local_adr==80) RDATA_80 <= WDATA;
	 if(local_adr==81) RDATA_81 <= WDATA;
	 if(local_adr==82) RDATA_82 <= WDATA;
	 if(local_adr==83) RDATA_83 <= WDATA;
	 if(local_adr==84) RDATA_84 <= WDATA;
	 if(local_adr==85) RDATA_85 <= WDATA;
	 if(local_adr==86) RDATA_86 <= WDATA;
	 if(local_adr==87) RDATA_87 <= WDATA;
	 if(local_adr==88) RDATA_88 <= WDATA;
	 if(local_adr==89) RDATA_89 <= WDATA;
	 if(local_adr==90) RDATA_90 <= WDATA;
	 if(local_adr==91) RDATA_91 <= WDATA;
	 if(local_adr==92) RDATA_92 <= WDATA;
	 if(local_adr==93) RDATA_93 <= WDATA;
	 if(local_adr==94) RDATA_94 <= WDATA;
	 if(local_adr==95) RDATA_95 <= WDATA;
	 if(local_adr==96) RDATA_96 <= WDATA;
	 if(local_adr==97) RDATA_97 <= WDATA;
	 if(local_adr==98) RDATA_98 <= WDATA;
	 if(local_adr==99) RDATA_99 <= WDATA;
	 if(local_adr==100) RDATA_100 <= WDATA;
	 if(local_adr==101) RDATA_101 <= WDATA;
	 if(local_adr==102) RDATA_102 <= WDATA;
	 if(local_adr==103) RDATA_103 <= WDATA;
	 if(local_adr==104) RDATA_104 <= WDATA;
	 if(local_adr==105) RDATA_105 <= WDATA;
	 if(local_adr==106) RDATA_106 <= WDATA;
	 if(local_adr==107) RDATA_107 <= WDATA;
	 if(local_adr==108) RDATA_108 <= WDATA;
	 if(local_adr==109) RDATA_109 <= WDATA;
	 if(local_adr==110) RDATA_110 <= WDATA;
	 if(local_adr==111) RDATA_111 <= WDATA;
	 if(local_adr==112) RDATA_112 <= WDATA;
	 if(local_adr==113) RDATA_113 <= WDATA;
	 if(local_adr==114) RDATA_114 <= WDATA;
	 if(local_adr==115) RDATA_115 <= WDATA;
	 if(local_adr==116) RDATA_116 <= WDATA;
	 if(local_adr==117) RDATA_117 <= WDATA;
	 if(local_adr==118) RDATA_118 <= WDATA;
	 if(local_adr==119) RDATA_119 <= WDATA;
	 if(local_adr==120) RDATA_120 <= WDATA;
	 if(local_adr==121) RDATA_121 <= WDATA;
	 if(local_adr==122) RDATA_122 <= WDATA;
	 if(local_adr==123) RDATA_123 <= WDATA;
	 if(local_adr==124) RDATA_124 <= WDATA;
	 if(local_adr==125) RDATA_125 <= WDATA;
	 if(local_adr==126) RDATA_126 <= WDATA;
	 if(local_adr==127) RDATA_127 <= WDATA;
	 if(local_adr==128) RDATA_128 <= WDATA;
	 if(local_adr==129) RDATA_129 <= WDATA;
	 if(local_adr==130) RDATA_130 <= WDATA;
	 if(local_adr==131) RDATA_131 <= WDATA;
	 if(local_adr==132) RDATA_132 <= WDATA;
	 if(local_adr==133) RDATA_133 <= WDATA;
	 if(local_adr==134) RDATA_134 <= WDATA;
	 if(local_adr==135) RDATA_135 <= WDATA;
	 if(local_adr==136) RDATA_136 <= WDATA;
	 if(local_adr==137) RDATA_137 <= WDATA;
	 if(local_adr==138) RDATA_138 <= WDATA;
	 if(local_adr==139) RDATA_139 <= WDATA;
	 if(local_adr==140) RDATA_140 <= WDATA;
	 if(local_adr==141) RDATA_141 <= WDATA;
	 if(local_adr==142) RDATA_142 <= WDATA;
	 if(local_adr==143) RDATA_143 <= WDATA;
	 if(local_adr==144) RDATA_144 <= WDATA;
	 if(local_adr==145) RDATA_145 <= WDATA;
	 if(local_adr==146) RDATA_146 <= WDATA;
	 if(local_adr==147) RDATA_147 <= WDATA;
	 if(local_adr==148) RDATA_148 <= WDATA;
	 if(local_adr==149) RDATA_149 <= WDATA;
	 if(local_adr==150) RDATA_150 <= WDATA;
	 if(local_adr==151) RDATA_151 <= WDATA;
	 if(local_adr==152) RDATA_152 <= WDATA;
	 if(local_adr==153) RDATA_153 <= WDATA;
	 if(local_adr==154) RDATA_154 <= WDATA;
	 if(local_adr==155) RDATA_155 <= WDATA;
	 if(local_adr==156) RDATA_156 <= WDATA;
	 if(local_adr==157) RDATA_157 <= WDATA;
	 if(local_adr==158) RDATA_158 <= WDATA;
	 if(local_adr==159) RDATA_159 <= WDATA;
	 if(local_adr==160) RDATA_160 <= WDATA;
	 if(local_adr==161) RDATA_161 <= WDATA;
	 if(local_adr==162) RDATA_162 <= WDATA;
	 if(local_adr==163) RDATA_163 <= WDATA;
	 if(local_adr==164) RDATA_164 <= WDATA;
	 if(local_adr==165) RDATA_165 <= WDATA;
	 if(local_adr==166) RDATA_166 <= WDATA;
	 if(local_adr==167) RDATA_167 <= WDATA;
	 if(local_adr==168) RDATA_168 <= WDATA;
	 if(local_adr==169) RDATA_169 <= WDATA;
	 if(local_adr==170) RDATA_170 <= WDATA;
	 if(local_adr==171) RDATA_171 <= WDATA;
	 if(local_adr==172) RDATA_172 <= WDATA;
	 if(local_adr==173) RDATA_173 <= WDATA;
	 if(local_adr==174) RDATA_174 <= WDATA;
	 if(local_adr==175) RDATA_175 <= WDATA;
	 if(local_adr==176) RDATA_176 <= WDATA;
	 if(local_adr==177) RDATA_177 <= WDATA;
	 if(local_adr==178) RDATA_178 <= WDATA;
	 if(local_adr==179) RDATA_179 <= WDATA;
	 if(local_adr==180) RDATA_180 <= WDATA;
	 if(local_adr==181) RDATA_181 <= WDATA;
	 if(local_adr==182) RDATA_182 <= WDATA;
	 if(local_adr==183) RDATA_183 <= WDATA;
	 if(local_adr==184) RDATA_184 <= WDATA;
	 if(local_adr==185) RDATA_185 <= WDATA;
	 if(local_adr==186) RDATA_186 <= WDATA;
	 if(local_adr==187) RDATA_187 <= WDATA;
	 if(local_adr==188) RDATA_188 <= WDATA;
	 if(local_adr==189) RDATA_189 <= WDATA;
	 if(local_adr==190) RDATA_190 <= WDATA;
	 if(local_adr==191) RDATA_191 <= WDATA;
	 if(local_adr==192) RDATA_192 <= WDATA;
	 if(local_adr==193) RDATA_193 <= WDATA;
	 if(local_adr==194) RDATA_194 <= WDATA;
	 if(local_adr==195) RDATA_195 <= WDATA;
	 if(local_adr==196) RDATA_196 <= WDATA;
	 if(local_adr==197) RDATA_197 <= WDATA;
	 if(local_adr==198) RDATA_198 <= WDATA;
	 if(local_adr==199) RDATA_199 <= WDATA;
	 if(local_adr==200) RDATA_200 <= WDATA;
	 if(local_adr==201) RDATA_201 <= WDATA;
	 if(local_adr==202) RDATA_202 <= WDATA;
	 if(local_adr==203) RDATA_203 <= WDATA;
	 if(local_adr==204) RDATA_204 <= WDATA;
	 if(local_adr==205) RDATA_205 <= WDATA;
	 if(local_adr==206) RDATA_206 <= WDATA;
	 if(local_adr==207) RDATA_207 <= WDATA;
	 if(local_adr==208) RDATA_208 <= WDATA;
	 if(local_adr==209) RDATA_209 <= WDATA;
	 if(local_adr==210) RDATA_210 <= WDATA;
	 if(local_adr==211) RDATA_211 <= WDATA;
	 if(local_adr==212) RDATA_212 <= WDATA;
	 if(local_adr==213) RDATA_213 <= WDATA;
	 if(local_adr==214) RDATA_214 <= WDATA;
	 if(local_adr==215) RDATA_215 <= WDATA;
	 if(local_adr==216) RDATA_216 <= WDATA;
	 if(local_adr==217) RDATA_217 <= WDATA;
	 if(local_adr==218) RDATA_218 <= WDATA;
	 if(local_adr==219) RDATA_219 <= WDATA;
	 if(local_adr==220) RDATA_220 <= WDATA;
	 if(local_adr==221) RDATA_221 <= WDATA;
	 if(local_adr==222) RDATA_222 <= WDATA;
	 if(local_adr==223) RDATA_223 <= WDATA;
	 if(local_adr==224) RDATA_224 <= WDATA;
	 if(local_adr==225) RDATA_225 <= WDATA;
	 if(local_adr==226) RDATA_226 <= WDATA;
	 if(local_adr==227) RDATA_227 <= WDATA;
	 if(local_adr==228) RDATA_228 <= WDATA;
	 if(local_adr==229) RDATA_229 <= WDATA;
	 if(local_adr==230) RDATA_230 <= WDATA;
	 if(local_adr==231) RDATA_231 <= WDATA;
	 if(local_adr==232) RDATA_232 <= WDATA;
	 if(local_adr==233) RDATA_233 <= WDATA;
	 if(local_adr==234) RDATA_234 <= WDATA;
	 if(local_adr==235) RDATA_235 <= WDATA;
	 if(local_adr==236) RDATA_236 <= WDATA;
	 if(local_adr==237) RDATA_237 <= WDATA;
	 if(local_adr==238) RDATA_238 <= WDATA;
	 if(local_adr==239) RDATA_239 <= WDATA;
	 if(local_adr==240) RDATA_240 <= WDATA;
	 if(local_adr==241) RDATA_241 <= WDATA;
	 if(local_adr==242) RDATA_242 <= WDATA;
	 if(local_adr==243) RDATA_243 <= WDATA;
	 if(local_adr==244) RDATA_244 <= WDATA;
	 if(local_adr==245) RDATA_245 <= WDATA;
	 if(local_adr==246) RDATA_246 <= WDATA;
	 if(local_adr==247) RDATA_247 <= WDATA;
	 if(local_adr==248) RDATA_248 <= WDATA;
	 if(local_adr==249) RDATA_249 <= WDATA;
	 if(local_adr==250) RDATA_250 <= WDATA;
	 if(local_adr==251) RDATA_251 <= WDATA;
	 if(local_adr==252) RDATA_252 <= WDATA;
	 if(local_adr==253) RDATA_253 <= WDATA;
	 if(local_adr==254) RDATA_254 <= WDATA;
	 if(local_adr==255) RDATA_255 <= WDATA;
	 if(local_adr==256) RDATA_256 <= WDATA;
	 if(local_adr==257) RDATA_257 <= WDATA;
	 if(local_adr==258) RDATA_258 <= WDATA;
	 if(local_adr==259) RDATA_259 <= WDATA;
	 if(local_adr==260) RDATA_260 <= WDATA;
	 if(local_adr==261) RDATA_261 <= WDATA;
	 if(local_adr==262) RDATA_262 <= WDATA;
	 if(local_adr==263) RDATA_263 <= WDATA;
	 if(local_adr==264) RDATA_264 <= WDATA;
	 if(local_adr==265) RDATA_265 <= WDATA;
	 if(local_adr==266) RDATA_266 <= WDATA;
	 if(local_adr==267) RDATA_267 <= WDATA;
	 if(local_adr==268) RDATA_268 <= WDATA;
	 if(local_adr==269) RDATA_269 <= WDATA;
	 if(local_adr==270) RDATA_270 <= WDATA;
	 if(local_adr==271) RDATA_271 <= WDATA;
	 if(local_adr==272) RDATA_272 <= WDATA;
	 if(local_adr==273) RDATA_273 <= WDATA;
	 if(local_adr==274) RDATA_274 <= WDATA;
	 if(local_adr==275) RDATA_275 <= WDATA;
	 if(local_adr==276) RDATA_276 <= WDATA;
	 if(local_adr==277) RDATA_277 <= WDATA;
	 if(local_adr==278) RDATA_278 <= WDATA;
	 if(local_adr==279) RDATA_279 <= WDATA;
	 if(local_adr==280) RDATA_280 <= WDATA;
	 if(local_adr==281) RDATA_281 <= WDATA;
	 if(local_adr==282) RDATA_282 <= WDATA;
	 if(local_adr==283) RDATA_283 <= WDATA;
	 if(local_adr==284) RDATA_284 <= WDATA;
	 if(local_adr==285) RDATA_285 <= WDATA;
	 if(local_adr==286) RDATA_286 <= WDATA;
	 if(local_adr==287) RDATA_287 <= WDATA;
	 if(local_adr==288) RDATA_288 <= WDATA;
	 if(local_adr==289) RDATA_289 <= WDATA;
	 if(local_adr==290) RDATA_290 <= WDATA;
	 if(local_adr==291) RDATA_291 <= WDATA;
	 if(local_adr==292) RDATA_292 <= WDATA;
	 if(local_adr==293) RDATA_293 <= WDATA;
	 if(local_adr==294) RDATA_294 <= WDATA;
	 if(local_adr==295) RDATA_295 <= WDATA;
	 if(local_adr==296) RDATA_296 <= WDATA;
	 if(local_adr==297) RDATA_297 <= WDATA;
	 if(local_adr==298) RDATA_298 <= WDATA;
	 if(local_adr==299) RDATA_299 <= WDATA;
	 if(local_adr==300) RDATA_300 <= WDATA;
	 if(local_adr==301) RDATA_301 <= WDATA;
	 if(local_adr==302) RDATA_302 <= WDATA;
	 if(local_adr==303) RDATA_303 <= WDATA;
	 if(local_adr==304) RDATA_304 <= WDATA;
	 if(local_adr==305) RDATA_305 <= WDATA;
	 if(local_adr==306) RDATA_306 <= WDATA;
	 if(local_adr==307) RDATA_307 <= WDATA;
	 if(local_adr==308) RDATA_308 <= WDATA;
	 if(local_adr==309) RDATA_309 <= WDATA;
	 if(local_adr==310) RDATA_310 <= WDATA;
	 if(local_adr==311) RDATA_311 <= WDATA;
	 if(local_adr==312) RDATA_312 <= WDATA;
	 if(local_adr==313) RDATA_313 <= WDATA;
	 if(local_adr==314) RDATA_314 <= WDATA;
	 if(local_adr==315) RDATA_315 <= WDATA;
	 if(local_adr==316) RDATA_316 <= WDATA;
	 if(local_adr==317) RDATA_317 <= WDATA;
	 if(local_adr==318) RDATA_318 <= WDATA;
	 if(local_adr==319) RDATA_319 <= WDATA;
	 if(local_adr==320) RDATA_320 <= WDATA;
	 if(local_adr==321) RDATA_321 <= WDATA;
	 if(local_adr==322) RDATA_322 <= WDATA;
	 if(local_adr==323) RDATA_323 <= WDATA;
	 if(local_adr==324) RDATA_324 <= WDATA;
	 if(local_adr==325) RDATA_325 <= WDATA;
	 if(local_adr==326) RDATA_326 <= WDATA;
	 if(local_adr==327) RDATA_327 <= WDATA;
	 if(local_adr==328) RDATA_328 <= WDATA;
	 if(local_adr==329) RDATA_329 <= WDATA;
	 if(local_adr==330) RDATA_330 <= WDATA;
	 if(local_adr==331) RDATA_331 <= WDATA;
	 if(local_adr==332) RDATA_332 <= WDATA;
	 if(local_adr==333) RDATA_333 <= WDATA;
	 if(local_adr==334) RDATA_334 <= WDATA;
	 if(local_adr==335) RDATA_335 <= WDATA;
	 if(local_adr==336) RDATA_336 <= WDATA;
	 if(local_adr==337) RDATA_337 <= WDATA;
	 if(local_adr==338) RDATA_338 <= WDATA;
	 if(local_adr==339) RDATA_339 <= WDATA;
	 if(local_adr==340) RDATA_340 <= WDATA;
	 if(local_adr==341) RDATA_341 <= WDATA;
	 if(local_adr==342) RDATA_342 <= WDATA;
	 if(local_adr==343) RDATA_343 <= WDATA;
	 if(local_adr==344) RDATA_344 <= WDATA;
	 if(local_adr==345) RDATA_345 <= WDATA;
	 if(local_adr==346) RDATA_346 <= WDATA;
	 if(local_adr==347) RDATA_347 <= WDATA;
	 if(local_adr==348) RDATA_348 <= WDATA;
	 if(local_adr==349) RDATA_349 <= WDATA;
	 if(local_adr==350) RDATA_350 <= WDATA;
	 if(local_adr==351) RDATA_351 <= WDATA;
	 if(local_adr==352) RDATA_352 <= WDATA;
	 if(local_adr==353) RDATA_353 <= WDATA;
	 if(local_adr==354) RDATA_354 <= WDATA;
	 if(local_adr==355) RDATA_355 <= WDATA;
	 if(local_adr==356) RDATA_356 <= WDATA;
	 if(local_adr==357) RDATA_357 <= WDATA;
	 if(local_adr==358) RDATA_358 <= WDATA;
	 if(local_adr==359) RDATA_359 <= WDATA;
	 if(local_adr==360) RDATA_360 <= WDATA;
	 if(local_adr==361) RDATA_361 <= WDATA;
	 if(local_adr==362) RDATA_362 <= WDATA;
	 if(local_adr==363) RDATA_363 <= WDATA;
	 if(local_adr==364) RDATA_364 <= WDATA;
	 if(local_adr==365) RDATA_365 <= WDATA;
	 if(local_adr==366) RDATA_366 <= WDATA;
	 if(local_adr==367) RDATA_367 <= WDATA;
	 if(local_adr==368) RDATA_368 <= WDATA;
	 if(local_adr==369) RDATA_369 <= WDATA;
	 if(local_adr==370) RDATA_370 <= WDATA;
	 if(local_adr==371) RDATA_371 <= WDATA;
	 if(local_adr==372) RDATA_372 <= WDATA;
	 if(local_adr==373) RDATA_373 <= WDATA;
	 if(local_adr==374) RDATA_374 <= WDATA;
	 if(local_adr==375) RDATA_375 <= WDATA;
	 if(local_adr==376) RDATA_376 <= WDATA;
	 if(local_adr==377) RDATA_377 <= WDATA;
	 if(local_adr==378) RDATA_378 <= WDATA;
	 if(local_adr==379) RDATA_379 <= WDATA;
	 if(local_adr==380) RDATA_380 <= WDATA;
	 if(local_adr==381) RDATA_381 <= WDATA;
	 if(local_adr==382) RDATA_382 <= WDATA;
	 if(local_adr==383) RDATA_383 <= WDATA;
	 if(local_adr==384) RDATA_384 <= WDATA;
	 if(local_adr==385) RDATA_385 <= WDATA;
	 if(local_adr==386) RDATA_386 <= WDATA;
	 if(local_adr==387) RDATA_387 <= WDATA;
	 if(local_adr==388) RDATA_388 <= WDATA;
	 if(local_adr==389) RDATA_389 <= WDATA;
	 if(local_adr==390) RDATA_390 <= WDATA;
	 if(local_adr==391) RDATA_391 <= WDATA;
	 if(local_adr==392) RDATA_392 <= WDATA;
	 if(local_adr==393) RDATA_393 <= WDATA;
	 if(local_adr==394) RDATA_394 <= WDATA;
	 if(local_adr==395) RDATA_395 <= WDATA;
	 if(local_adr==396) RDATA_396 <= WDATA;
	 if(local_adr==397) RDATA_397 <= WDATA;
	 if(local_adr==398) RDATA_398 <= WDATA;
	 if(local_adr==399) RDATA_399 <= WDATA;
	 if(local_adr==400) RDATA_400 <= WDATA;
	 if(local_adr==401) RDATA_401 <= WDATA;
	 if(local_adr==402) RDATA_402 <= WDATA;
	 if(local_adr==403) RDATA_403 <= WDATA;
	 if(local_adr==404) RDATA_404 <= WDATA;
	 if(local_adr==405) RDATA_405 <= WDATA;
	 if(local_adr==406) RDATA_406 <= WDATA;
	 if(local_adr==407) RDATA_407 <= WDATA;
	 if(local_adr==408) RDATA_408 <= WDATA;
	 if(local_adr==409) RDATA_409 <= WDATA;
	 if(local_adr==410) RDATA_410 <= WDATA;
	 if(local_adr==411) RDATA_411 <= WDATA;
	 if(local_adr==412) RDATA_412 <= WDATA;
	 if(local_adr==413) RDATA_413 <= WDATA;
	 if(local_adr==414) RDATA_414 <= WDATA;
	 if(local_adr==415) RDATA_415 <= WDATA;
	 if(local_adr==416) RDATA_416 <= WDATA;
	 if(local_adr==417) RDATA_417 <= WDATA;
	 if(local_adr==418) RDATA_418 <= WDATA;
	 if(local_adr==419) RDATA_419 <= WDATA;
	 if(local_adr==420) RDATA_420 <= WDATA;
	 if(local_adr==421) RDATA_421 <= WDATA;
	 if(local_adr==422) RDATA_422 <= WDATA;
	 if(local_adr==423) RDATA_423 <= WDATA;
	 if(local_adr==424) RDATA_424 <= WDATA;
	 if(local_adr==425) RDATA_425 <= WDATA;
	 if(local_adr==426) RDATA_426 <= WDATA;
	 if(local_adr==427) RDATA_427 <= WDATA;
	 if(local_adr==428) RDATA_428 <= WDATA;
	 if(local_adr==429) RDATA_429 <= WDATA;
	 if(local_adr==430) RDATA_430 <= WDATA;
	 if(local_adr==431) RDATA_431 <= WDATA;
	 if(local_adr==432) RDATA_432 <= WDATA;
	 if(local_adr==433) RDATA_433 <= WDATA;
	 if(local_adr==434) RDATA_434 <= WDATA;
	 if(local_adr==435) RDATA_435 <= WDATA;
	 if(local_adr==436) RDATA_436 <= WDATA;
	 if(local_adr==437) RDATA_437 <= WDATA;
	 if(local_adr==438) RDATA_438 <= WDATA;
	 if(local_adr==439) RDATA_439 <= WDATA;
	 if(local_adr==440) RDATA_440 <= WDATA;
	 if(local_adr==441) RDATA_441 <= WDATA;
	 if(local_adr==442) RDATA_442 <= WDATA;
	 if(local_adr==443) RDATA_443 <= WDATA;
	 if(local_adr==444) RDATA_444 <= WDATA;
	 if(local_adr==445) RDATA_445 <= WDATA;
	 if(local_adr==446) RDATA_446 <= WDATA;
	 if(local_adr==447) RDATA_447 <= WDATA;
	 if(local_adr==448) RDATA_448 <= WDATA;
	 if(local_adr==449) RDATA_449 <= WDATA;
	 if(local_adr==450) RDATA_450 <= WDATA;
	 if(local_adr==451) RDATA_451 <= WDATA;
	 if(local_adr==452) RDATA_452 <= WDATA;
	 if(local_adr==453) RDATA_453 <= WDATA;
	 if(local_adr==454) RDATA_454 <= WDATA;
	 if(local_adr==455) RDATA_455 <= WDATA;
	 if(local_adr==456) RDATA_456 <= WDATA;
	 if(local_adr==457) RDATA_457 <= WDATA;
	 if(local_adr==458) RDATA_458 <= WDATA;
	 if(local_adr==459) RDATA_459 <= WDATA;
	 if(local_adr==460) RDATA_460 <= WDATA;
	 if(local_adr==461) RDATA_461 <= WDATA;
	 if(local_adr==462) RDATA_462 <= WDATA;
	 if(local_adr==463) RDATA_463 <= WDATA;
	 if(local_adr==464) RDATA_464 <= WDATA;
	 if(local_adr==465) RDATA_465 <= WDATA;
	 if(local_adr==466) RDATA_466 <= WDATA;
	 if(local_adr==467) RDATA_467 <= WDATA;
	 if(local_adr==468) RDATA_468 <= WDATA;
	 if(local_adr==469) RDATA_469 <= WDATA;
	 if(local_adr==470) RDATA_470 <= WDATA;
	 if(local_adr==471) RDATA_471 <= WDATA;
	 if(local_adr==472) RDATA_472 <= WDATA;
	 if(local_adr==473) RDATA_473 <= WDATA;
	 if(local_adr==474) RDATA_474 <= WDATA;
	 if(local_adr==475) RDATA_475 <= WDATA;
	 if(local_adr==476) RDATA_476 <= WDATA;
	 if(local_adr==477) RDATA_477 <= WDATA;
	 if(local_adr==478) RDATA_478 <= WDATA;
	 if(local_adr==479) RDATA_479 <= WDATA;
	 if(local_adr==480) RDATA_480 <= WDATA;
	 if(local_adr==481) RDATA_481 <= WDATA;
	 if(local_adr==482) RDATA_482 <= WDATA;
	 if(local_adr==483) RDATA_483 <= WDATA;
	 if(local_adr==484) RDATA_484 <= WDATA;
	 if(local_adr==485) RDATA_485 <= WDATA;
	 if(local_adr==486) RDATA_486 <= WDATA;
	 if(local_adr==487) RDATA_487 <= WDATA;
	 if(local_adr==488) RDATA_488 <= WDATA;
	 if(local_adr==489) RDATA_489 <= WDATA;
	 if(local_adr==490) RDATA_490 <= WDATA;
	 if(local_adr==491) RDATA_491 <= WDATA;
	 if(local_adr==492) RDATA_492 <= WDATA;
	 if(local_adr==493) RDATA_493 <= WDATA;
	 if(local_adr==494) RDATA_494 <= WDATA;
	 if(local_adr==495) RDATA_495 <= WDATA;
	 if(local_adr==496) RDATA_496 <= WDATA;
	 if(local_adr==497) RDATA_497 <= WDATA;
	 if(local_adr==498) RDATA_498 <= WDATA;
	 if(local_adr==499) RDATA_499 <= WDATA;
	 if(local_adr==500) RDATA_500 <= WDATA;
	 if(local_adr==501) RDATA_501 <= WDATA;
	 if(local_adr==502) RDATA_502 <= WDATA;
	 if(local_adr==503) RDATA_503 <= WDATA;
	 if(local_adr==504) RDATA_504 <= WDATA;
	 if(local_adr==505) RDATA_505 <= WDATA;
	 if(local_adr==506) RDATA_506 <= WDATA;
	 if(local_adr==507) RDATA_507 <= WDATA;
	 if(local_adr==508) RDATA_508 <= WDATA;
	 if(local_adr==509) RDATA_509 <= WDATA;
	 if(local_adr==510) RDATA_510 <= WDATA;
	 if(local_adr==511) RDATA_511 <= WDATA;
	 if(local_adr==512) RDATA_512 <= WDATA;
	 if(local_adr==513) RDATA_513 <= WDATA;
	 if(local_adr==514) RDATA_514 <= WDATA;
	 if(local_adr==515) RDATA_515 <= WDATA;
	 if(local_adr==516) RDATA_516 <= WDATA;
	 if(local_adr==517) RDATA_517 <= WDATA;
	 if(local_adr==518) RDATA_518 <= WDATA;
	 if(local_adr==519) RDATA_519 <= WDATA;
	 if(local_adr==520) RDATA_520 <= WDATA;
	 if(local_adr==521) RDATA_521 <= WDATA;
	 if(local_adr==522) RDATA_522 <= WDATA;
	 if(local_adr==523) RDATA_523 <= WDATA;
	 if(local_adr==524) RDATA_524 <= WDATA;
	 if(local_adr==525) RDATA_525 <= WDATA;
	 if(local_adr==526) RDATA_526 <= WDATA;
	 if(local_adr==527) RDATA_527 <= WDATA;
	 if(local_adr==528) RDATA_528 <= WDATA;
	 if(local_adr==529) RDATA_529 <= WDATA;
	 if(local_adr==530) RDATA_530 <= WDATA;
	 if(local_adr==531) RDATA_531 <= WDATA;
	 if(local_adr==532) RDATA_532 <= WDATA;
	 if(local_adr==533) RDATA_533 <= WDATA;
	 if(local_adr==534) RDATA_534 <= WDATA;
	 if(local_adr==535) RDATA_535 <= WDATA;
	 if(local_adr==536) RDATA_536 <= WDATA;
	 if(local_adr==537) RDATA_537 <= WDATA;
	 if(local_adr==538) RDATA_538 <= WDATA;
	 if(local_adr==539) RDATA_539 <= WDATA;
	 if(local_adr==540) RDATA_540 <= WDATA;
	 if(local_adr==541) RDATA_541 <= WDATA;
	 if(local_adr==542) RDATA_542 <= WDATA;
	 if(local_adr==543) RDATA_543 <= WDATA;
	 if(local_adr==544) RDATA_544 <= WDATA;
	 if(local_adr==545) RDATA_545 <= WDATA;
	 if(local_adr==546) RDATA_546 <= WDATA;
	 if(local_adr==547) RDATA_547 <= WDATA;
	 if(local_adr==548) RDATA_548 <= WDATA;
	 if(local_adr==549) RDATA_549 <= WDATA;
	 if(local_adr==550) RDATA_550 <= WDATA;
	 if(local_adr==551) RDATA_551 <= WDATA;
	 if(local_adr==552) RDATA_552 <= WDATA;
	 if(local_adr==553) RDATA_553 <= WDATA;
	 if(local_adr==554) RDATA_554 <= WDATA;
	 if(local_adr==555) RDATA_555 <= WDATA;
	 if(local_adr==556) RDATA_556 <= WDATA;
	 if(local_adr==557) RDATA_557 <= WDATA;
	 if(local_adr==558) RDATA_558 <= WDATA;
	 if(local_adr==559) RDATA_559 <= WDATA;
	 if(local_adr==560) RDATA_560 <= WDATA;
	 if(local_adr==561) RDATA_561 <= WDATA;
	 if(local_adr==562) RDATA_562 <= WDATA;
	 if(local_adr==563) RDATA_563 <= WDATA;
	 if(local_adr==564) RDATA_564 <= WDATA;
	 if(local_adr==565) RDATA_565 <= WDATA;
	 if(local_adr==566) RDATA_566 <= WDATA;
	 if(local_adr==567) RDATA_567 <= WDATA;
	 if(local_adr==568) RDATA_568 <= WDATA;
	 if(local_adr==569) RDATA_569 <= WDATA;
	 if(local_adr==570) RDATA_570 <= WDATA;
	 if(local_adr==571) RDATA_571 <= WDATA;
	 if(local_adr==572) RDATA_572 <= WDATA;
	 if(local_adr==573) RDATA_573 <= WDATA;
	 if(local_adr==574) RDATA_574 <= WDATA;
	 if(local_adr==575) RDATA_575 <= WDATA;
	 if(local_adr==576) RDATA_576 <= WDATA;
	 if(local_adr==577) RDATA_577 <= WDATA;
	 if(local_adr==578) RDATA_578 <= WDATA;
	 if(local_adr==579) RDATA_579 <= WDATA;
	 if(local_adr==580) RDATA_580 <= WDATA;
	 if(local_adr==581) RDATA_581 <= WDATA;
	 if(local_adr==582) RDATA_582 <= WDATA;
	 if(local_adr==583) RDATA_583 <= WDATA;
	 if(local_adr==584) RDATA_584 <= WDATA;
	 if(local_adr==585) RDATA_585 <= WDATA;
	 if(local_adr==586) RDATA_586 <= WDATA;
	 if(local_adr==587) RDATA_587 <= WDATA;
	 if(local_adr==588) RDATA_588 <= WDATA;
	 if(local_adr==589) RDATA_589 <= WDATA;
	 if(local_adr==590) RDATA_590 <= WDATA;
	 if(local_adr==591) RDATA_591 <= WDATA;
	 if(local_adr==592) RDATA_592 <= WDATA;
	 if(local_adr==593) RDATA_593 <= WDATA;
	 if(local_adr==594) RDATA_594 <= WDATA;
	 if(local_adr==595) RDATA_595 <= WDATA;
	 if(local_adr==596) RDATA_596 <= WDATA;
	 if(local_adr==597) RDATA_597 <= WDATA;
	 if(local_adr==598) RDATA_598 <= WDATA;
	 if(local_adr==599) RDATA_599 <= WDATA;
	 if(local_adr==600) RDATA_600 <= WDATA;
	 if(local_adr==601) RDATA_601 <= WDATA;
	 if(local_adr==602) RDATA_602 <= WDATA;
	 if(local_adr==603) RDATA_603 <= WDATA;
	 if(local_adr==604) RDATA_604 <= WDATA;
	 if(local_adr==605) RDATA_605 <= WDATA;
	 if(local_adr==606) RDATA_606 <= WDATA;
	 if(local_adr==607) RDATA_607 <= WDATA;
	 if(local_adr==608) RDATA_608 <= WDATA;
	 if(local_adr==609) RDATA_609 <= WDATA;
	 if(local_adr==610) RDATA_610 <= WDATA;
	 if(local_adr==611) RDATA_611 <= WDATA;
	 if(local_adr==612) RDATA_612 <= WDATA;
	 if(local_adr==613) RDATA_613 <= WDATA;
	 if(local_adr==614) RDATA_614 <= WDATA;
	 if(local_adr==615) RDATA_615 <= WDATA;
	 if(local_adr==616) RDATA_616 <= WDATA;
	 if(local_adr==617) RDATA_617 <= WDATA;
	 if(local_adr==618) RDATA_618 <= WDATA;
	 if(local_adr==619) RDATA_619 <= WDATA;
	 if(local_adr==620) RDATA_620 <= WDATA;
	 if(local_adr==621) RDATA_621 <= WDATA;
	 if(local_adr==622) RDATA_622 <= WDATA;
	 if(local_adr==623) RDATA_623 <= WDATA;
	 if(local_adr==624) RDATA_624 <= WDATA;
	 if(local_adr==625) RDATA_625 <= WDATA;
	 if(local_adr==626) RDATA_626 <= WDATA;
	 if(local_adr==627) RDATA_627 <= WDATA;
	 if(local_adr==628) RDATA_628 <= WDATA;
	 if(local_adr==629) RDATA_629 <= WDATA;
	 if(local_adr==630) RDATA_630 <= WDATA;
	 if(local_adr==631) RDATA_631 <= WDATA;
	 if(local_adr==632) RDATA_632 <= WDATA;
	 if(local_adr==633) RDATA_633 <= WDATA;
	 if(local_adr==634) RDATA_634 <= WDATA;
	 if(local_adr==635) RDATA_635 <= WDATA;
	 if(local_adr==636) RDATA_636 <= WDATA;
	 if(local_adr==637) RDATA_637 <= WDATA;
	 if(local_adr==638) RDATA_638 <= WDATA;
	 if(local_adr==639) RDATA_639 <= WDATA;
	 if(local_adr==640) RDATA_640 <= WDATA;
	 if(local_adr==641) RDATA_641 <= WDATA;
	 if(local_adr==642) RDATA_642 <= WDATA;
	 if(local_adr==643) RDATA_643 <= WDATA;
	 if(local_adr==644) RDATA_644 <= WDATA;
	 if(local_adr==645) RDATA_645 <= WDATA;
	 if(local_adr==646) RDATA_646 <= WDATA;
	 if(local_adr==647) RDATA_647 <= WDATA;
	 if(local_adr==648) RDATA_648 <= WDATA;
	 if(local_adr==649) RDATA_649 <= WDATA;
	 if(local_adr==650) RDATA_650 <= WDATA;
	 if(local_adr==651) RDATA_651 <= WDATA;
	 if(local_adr==652) RDATA_652 <= WDATA;
	 if(local_adr==653) RDATA_653 <= WDATA;
	 if(local_adr==654) RDATA_654 <= WDATA;
	 if(local_adr==655) RDATA_655 <= WDATA;
	 if(local_adr==656) RDATA_656 <= WDATA;
	 if(local_adr==657) RDATA_657 <= WDATA;
	 if(local_adr==658) RDATA_658 <= WDATA;
	 if(local_adr==659) RDATA_659 <= WDATA;
	 if(local_adr==660) RDATA_660 <= WDATA;
	 if(local_adr==661) RDATA_661 <= WDATA;
	 if(local_adr==662) RDATA_662 <= WDATA;
	 if(local_adr==663) RDATA_663 <= WDATA;
	 if(local_adr==664) RDATA_664 <= WDATA;
	 if(local_adr==665) RDATA_665 <= WDATA;
	 if(local_adr==666) RDATA_666 <= WDATA;
	 if(local_adr==667) RDATA_667 <= WDATA;
	 if(local_adr==668) RDATA_668 <= WDATA;
	 if(local_adr==669) RDATA_669 <= WDATA;
	 if(local_adr==670) RDATA_670 <= WDATA;
	 if(local_adr==671) RDATA_671 <= WDATA;
	 if(local_adr==672) RDATA_672 <= WDATA;
	 if(local_adr==673) RDATA_673 <= WDATA;
	 if(local_adr==674) RDATA_674 <= WDATA;
	 if(local_adr==675) RDATA_675 <= WDATA;
	 if(local_adr==676) RDATA_676 <= WDATA;
	 if(local_adr==677) RDATA_677 <= WDATA;
	 if(local_adr==678) RDATA_678 <= WDATA;
	 if(local_adr==679) RDATA_679 <= WDATA;
	 if(local_adr==680) RDATA_680 <= WDATA;
	 if(local_adr==681) RDATA_681 <= WDATA;
	 if(local_adr==682) RDATA_682 <= WDATA;
	 if(local_adr==683) RDATA_683 <= WDATA;
	 if(local_adr==684) RDATA_684 <= WDATA;
	 if(local_adr==685) RDATA_685 <= WDATA;
	 if(local_adr==686) RDATA_686 <= WDATA;
	 if(local_adr==687) RDATA_687 <= WDATA;
	 if(local_adr==688) RDATA_688 <= WDATA;
	 if(local_adr==689) RDATA_689 <= WDATA;
	 if(local_adr==690) RDATA_690 <= WDATA;
	 if(local_adr==691) RDATA_691 <= WDATA;
	 if(local_adr==692) RDATA_692 <= WDATA;
	 if(local_adr==693) RDATA_693 <= WDATA;
	 if(local_adr==694) RDATA_694 <= WDATA;
	 if(local_adr==695) RDATA_695 <= WDATA;
	 if(local_adr==696) RDATA_696 <= WDATA;
	 if(local_adr==697) RDATA_697 <= WDATA;
	 if(local_adr==698) RDATA_698 <= WDATA;
	 if(local_adr==699) RDATA_699 <= WDATA;
	 if(local_adr==700) RDATA_700 <= WDATA;
	 if(local_adr==701) RDATA_701 <= WDATA;
	 if(local_adr==702) RDATA_702 <= WDATA;
	 if(local_adr==703) RDATA_703 <= WDATA;
	 if(local_adr==704) RDATA_704 <= WDATA;
	 if(local_adr==705) RDATA_705 <= WDATA;
	 if(local_adr==706) RDATA_706 <= WDATA;
	 if(local_adr==707) RDATA_707 <= WDATA;
	 if(local_adr==708) RDATA_708 <= WDATA;
	 if(local_adr==709) RDATA_709 <= WDATA;
	 if(local_adr==710) RDATA_710 <= WDATA;
	 if(local_adr==711) RDATA_711 <= WDATA;
	 if(local_adr==712) RDATA_712 <= WDATA;
	 if(local_adr==713) RDATA_713 <= WDATA;
	 if(local_adr==714) RDATA_714 <= WDATA;
	 if(local_adr==715) RDATA_715 <= WDATA;
	 if(local_adr==716) RDATA_716 <= WDATA;
	 if(local_adr==717) RDATA_717 <= WDATA;
	 if(local_adr==718) RDATA_718 <= WDATA;
	 if(local_adr==719) RDATA_719 <= WDATA;
	 if(local_adr==720) RDATA_720 <= WDATA;
	 if(local_adr==721) RDATA_721 <= WDATA;
	 if(local_adr==722) RDATA_722 <= WDATA;
	 if(local_adr==723) RDATA_723 <= WDATA;
	 if(local_adr==724) RDATA_724 <= WDATA;
	 if(local_adr==725) RDATA_725 <= WDATA;
	 if(local_adr==726) RDATA_726 <= WDATA;
	 if(local_adr==727) RDATA_727 <= WDATA;
	 if(local_adr==728) RDATA_728 <= WDATA;
	 if(local_adr==729) RDATA_729 <= WDATA;
	 if(local_adr==730) RDATA_730 <= WDATA;
	 if(local_adr==731) RDATA_731 <= WDATA;
	 if(local_adr==732) RDATA_732 <= WDATA;
	 if(local_adr==733) RDATA_733 <= WDATA;
	 if(local_adr==734) RDATA_734 <= WDATA;
	 if(local_adr==735) RDATA_735 <= WDATA;
	 if(local_adr==736) RDATA_736 <= WDATA;
	 if(local_adr==737) RDATA_737 <= WDATA;
	 if(local_adr==738) RDATA_738 <= WDATA;
	 if(local_adr==739) RDATA_739 <= WDATA;
	 if(local_adr==740) RDATA_740 <= WDATA;
	 if(local_adr==741) RDATA_741 <= WDATA;
	 if(local_adr==742) RDATA_742 <= WDATA;
	 if(local_adr==743) RDATA_743 <= WDATA;
	 if(local_adr==744) RDATA_744 <= WDATA;
	 if(local_adr==745) RDATA_745 <= WDATA;
	 if(local_adr==746) RDATA_746 <= WDATA;
	 if(local_adr==747) RDATA_747 <= WDATA;
	 if(local_adr==748) RDATA_748 <= WDATA;
	 if(local_adr==749) RDATA_749 <= WDATA;
	 if(local_adr==750) RDATA_750 <= WDATA;
	 if(local_adr==751) RDATA_751 <= WDATA;
	 if(local_adr==752) RDATA_752 <= WDATA;
	 if(local_adr==753) RDATA_753 <= WDATA;
	 if(local_adr==754) RDATA_754 <= WDATA;
	 if(local_adr==755) RDATA_755 <= WDATA;
	 if(local_adr==756) RDATA_756 <= WDATA;
	 if(local_adr==757) RDATA_757 <= WDATA;
	 if(local_adr==758) RDATA_758 <= WDATA;
	 if(local_adr==759) RDATA_759 <= WDATA;
	 if(local_adr==760) RDATA_760 <= WDATA;
	 if(local_adr==761) RDATA_761 <= WDATA;
	 if(local_adr==762) RDATA_762 <= WDATA;
	 if(local_adr==763) RDATA_763 <= WDATA;
	 if(local_adr==764) RDATA_764 <= WDATA;
	 if(local_adr==765) RDATA_765 <= WDATA;
	 if(local_adr==766) RDATA_766 <= WDATA;
	 if(local_adr==767) RDATA_767 <= WDATA;
	 if(local_adr==768) RDATA_768 <= WDATA;
	 if(local_adr==769) RDATA_769 <= WDATA;
	 if(local_adr==770) RDATA_770 <= WDATA;
	 if(local_adr==771) RDATA_771 <= WDATA;
	 if(local_adr==772) RDATA_772 <= WDATA;
	 if(local_adr==773) RDATA_773 <= WDATA;
	 if(local_adr==774) RDATA_774 <= WDATA;
	 if(local_adr==775) RDATA_775 <= WDATA;
	 if(local_adr==776) RDATA_776 <= WDATA;
	 if(local_adr==777) RDATA_777 <= WDATA;
	 if(local_adr==778) RDATA_778 <= WDATA;
	 if(local_adr==779) RDATA_779 <= WDATA;
	 if(local_adr==780) RDATA_780 <= WDATA;
	 if(local_adr==781) RDATA_781 <= WDATA;
	 if(local_adr==782) RDATA_782 <= WDATA;
	 if(local_adr==783) RDATA_783 <= WDATA;
      end
   end // always @ (posedge CLK)
   
   assign RDATA[7:0] = RDATA_00;
   assign RDATA[15:8] = RDATA_01;
   assign RDATA[23:16] = RDATA_02;
   assign RDATA[31:24] = RDATA_03;
   assign RDATA[39:32] = RDATA_04;
   assign RDATA[47:40] = RDATA_05;
   assign RDATA[55:48] = RDATA_06;
   assign RDATA[63:56] = RDATA_07;
   assign RDATA[71:64] = RDATA_08;
   assign RDATA[79:72] = RDATA_09;
   assign RDATA[87:80] = RDATA_10;
   assign RDATA[95:88] = RDATA_11;
   assign RDATA[103:96] = RDATA_12;
   assign RDATA[111:104] = RDATA_13;
   assign RDATA[119:112] = RDATA_14;
   assign RDATA[127:120] = RDATA_15;
   assign RDATA[135:128] = RDATA_16;
   assign RDATA[143:136] = RDATA_17;
   assign RDATA[151:144] = RDATA_18;
   assign RDATA[159:152] = RDATA_19;
   assign RDATA[167:160] = RDATA_20;
   assign RDATA[175:168] = RDATA_21;
   assign RDATA[183:176] = RDATA_22;
   assign RDATA[191:184] = RDATA_23;
   assign RDATA[199:192] = RDATA_24;
   assign RDATA[207:200] = RDATA_25;
   assign RDATA[215:208] = RDATA_26;
   assign RDATA[223:216] = RDATA_27;
   assign RDATA[231:224] = RDATA_28;
   assign RDATA[239:232] = RDATA_29;
   assign RDATA[247:240] = RDATA_30;
   assign RDATA[255:248] = RDATA_31;
   assign RDATA[263:256] = RDATA_32;
   assign RDATA[271:264] = RDATA_33;
   assign RDATA[279:272] = RDATA_34;
   assign RDATA[287:280] = RDATA_35;
   assign RDATA[295:288] = RDATA_36;
   assign RDATA[303:296] = RDATA_37;
   assign RDATA[311:304] = RDATA_38;
   assign RDATA[319:312] = RDATA_39;
   assign RDATA[327:320] = RDATA_40;
   assign RDATA[335:328] = RDATA_41;
   assign RDATA[343:336] = RDATA_42;
   assign RDATA[351:344] = RDATA_43;
   assign RDATA[359:352] = RDATA_44;
   assign RDATA[367:360] = RDATA_45;
   assign RDATA[375:368] = RDATA_46;
   assign RDATA[383:376] = RDATA_47;
   assign RDATA[391:384] = RDATA_48;
   assign RDATA[399:392] = RDATA_49;
   assign RDATA[407:400] = RDATA_50;
   assign RDATA[415:408] = RDATA_51;
   assign RDATA[423:416] = RDATA_52;
   assign RDATA[431:424] = RDATA_53;
   assign RDATA[439:432] = RDATA_54;
   assign RDATA[447:440] = RDATA_55;
   assign RDATA[455:448] = RDATA_56;
   assign RDATA[463:456] = RDATA_57;
   assign RDATA[471:464] = RDATA_58;
   assign RDATA[479:472] = RDATA_59;
   assign RDATA[487:480] = RDATA_60;
   assign RDATA[495:488] = RDATA_61;
   assign RDATA[503:496] = RDATA_62;
   assign RDATA[511:504] = RDATA_63;
   assign RDATA[519:512] = RDATA_64;
   assign RDATA[527:520] = RDATA_65;
   assign RDATA[535:528] = RDATA_66;
   assign RDATA[543:536] = RDATA_67;
   assign RDATA[551:544] = RDATA_68;
   assign RDATA[559:552] = RDATA_69;
   assign RDATA[567:560] = RDATA_70;
   assign RDATA[575:568] = RDATA_71;
   assign RDATA[583:576] = RDATA_72;
   assign RDATA[591:584] = RDATA_73;
   assign RDATA[599:592] = RDATA_74;
   assign RDATA[607:600] = RDATA_75;
   assign RDATA[615:608] = RDATA_76;
   assign RDATA[623:616] = RDATA_77;
   assign RDATA[631:624] = RDATA_78;
   assign RDATA[639:632] = RDATA_79;
   assign RDATA[647:640] = RDATA_80;
   assign RDATA[655:648] = RDATA_81;
   assign RDATA[663:656] = RDATA_82;
   assign RDATA[671:664] = RDATA_83;
   assign RDATA[679:672] = RDATA_84;
   assign RDATA[687:680] = RDATA_85;
   assign RDATA[695:688] = RDATA_86;
   assign RDATA[703:696] = RDATA_87;
   assign RDATA[711:704] = RDATA_88;
   assign RDATA[719:712] = RDATA_89;
   assign RDATA[727:720] = RDATA_90;
   assign RDATA[735:728] = RDATA_91;
   assign RDATA[743:736] = RDATA_92;
   assign RDATA[751:744] = RDATA_93;
   assign RDATA[759:752] = RDATA_94;
   assign RDATA[767:760] = RDATA_95;
   assign RDATA[775:768] = RDATA_96;
   assign RDATA[783:776] = RDATA_97;
   assign RDATA[791:784] = RDATA_98;
   assign RDATA[799:792] = RDATA_99;
   assign RDATA[807:800] = RDATA_100;
   assign RDATA[815:808] = RDATA_101;
   assign RDATA[823:816] = RDATA_102;
   assign RDATA[831:824] = RDATA_103;
   assign RDATA[839:832] = RDATA_104;
   assign RDATA[847:840] = RDATA_105;
   assign RDATA[855:848] = RDATA_106;
   assign RDATA[863:856] = RDATA_107;
   assign RDATA[871:864] = RDATA_108;
   assign RDATA[879:872] = RDATA_109;
   assign RDATA[887:880] = RDATA_110;
   assign RDATA[895:888] = RDATA_111;
   assign RDATA[903:896] = RDATA_112;
   assign RDATA[911:904] = RDATA_113;
   assign RDATA[919:912] = RDATA_114;
   assign RDATA[927:920] = RDATA_115;
   assign RDATA[935:928] = RDATA_116;
   assign RDATA[943:936] = RDATA_117;
   assign RDATA[951:944] = RDATA_118;
   assign RDATA[959:952] = RDATA_119;
   assign RDATA[967:960] = RDATA_120;
   assign RDATA[975:968] = RDATA_121;
   assign RDATA[983:976] = RDATA_122;
   assign RDATA[991:984] = RDATA_123;
   assign RDATA[999:992] = RDATA_124;
   assign RDATA[1007:1000] = RDATA_125;
   assign RDATA[1015:1008] = RDATA_126;
   assign RDATA[1023:1016] = RDATA_127;
   assign RDATA[1031:1024] = RDATA_128;
   assign RDATA[1039:1032] = RDATA_129;
   assign RDATA[1047:1040] = RDATA_130;
   assign RDATA[1055:1048] = RDATA_131;
   assign RDATA[1063:1056] = RDATA_132;
   assign RDATA[1071:1064] = RDATA_133;
   assign RDATA[1079:1072] = RDATA_134;
   assign RDATA[1087:1080] = RDATA_135;
   assign RDATA[1095:1088] = RDATA_136;
   assign RDATA[1103:1096] = RDATA_137;
   assign RDATA[1111:1104] = RDATA_138;
   assign RDATA[1119:1112] = RDATA_139;
   assign RDATA[1127:1120] = RDATA_140;
   assign RDATA[1135:1128] = RDATA_141;
   assign RDATA[1143:1136] = RDATA_142;
   assign RDATA[1151:1144] = RDATA_143;
   assign RDATA[1159:1152] = RDATA_144;
   assign RDATA[1167:1160] = RDATA_145;
   assign RDATA[1175:1168] = RDATA_146;
   assign RDATA[1183:1176] = RDATA_147;
   assign RDATA[1191:1184] = RDATA_148;
   assign RDATA[1199:1192] = RDATA_149;
   assign RDATA[1207:1200] = RDATA_150;
   assign RDATA[1215:1208] = RDATA_151;
   assign RDATA[1223:1216] = RDATA_152;
   assign RDATA[1231:1224] = RDATA_153;
   assign RDATA[1239:1232] = RDATA_154;
   assign RDATA[1247:1240] = RDATA_155;
   assign RDATA[1255:1248] = RDATA_156;
   assign RDATA[1263:1256] = RDATA_157;
   assign RDATA[1271:1264] = RDATA_158;
   assign RDATA[1279:1272] = RDATA_159;
   assign RDATA[1287:1280] = RDATA_160;
   assign RDATA[1295:1288] = RDATA_161;
   assign RDATA[1303:1296] = RDATA_162;
   assign RDATA[1311:1304] = RDATA_163;
   assign RDATA[1319:1312] = RDATA_164;
   assign RDATA[1327:1320] = RDATA_165;
   assign RDATA[1335:1328] = RDATA_166;
   assign RDATA[1343:1336] = RDATA_167;
   assign RDATA[1351:1344] = RDATA_168;
   assign RDATA[1359:1352] = RDATA_169;
   assign RDATA[1367:1360] = RDATA_170;
   assign RDATA[1375:1368] = RDATA_171;
   assign RDATA[1383:1376] = RDATA_172;
   assign RDATA[1391:1384] = RDATA_173;
   assign RDATA[1399:1392] = RDATA_174;
   assign RDATA[1407:1400] = RDATA_175;
   assign RDATA[1415:1408] = RDATA_176;
   assign RDATA[1423:1416] = RDATA_177;
   assign RDATA[1431:1424] = RDATA_178;
   assign RDATA[1439:1432] = RDATA_179;
   assign RDATA[1447:1440] = RDATA_180;
   assign RDATA[1455:1448] = RDATA_181;
   assign RDATA[1463:1456] = RDATA_182;
   assign RDATA[1471:1464] = RDATA_183;
   assign RDATA[1479:1472] = RDATA_184;
   assign RDATA[1487:1480] = RDATA_185;
   assign RDATA[1495:1488] = RDATA_186;
   assign RDATA[1503:1496] = RDATA_187;
   assign RDATA[1511:1504] = RDATA_188;
   assign RDATA[1519:1512] = RDATA_189;
   assign RDATA[1527:1520] = RDATA_190;
   assign RDATA[1535:1528] = RDATA_191;
   assign RDATA[1543:1536] = RDATA_192;
   assign RDATA[1551:1544] = RDATA_193;
   assign RDATA[1559:1552] = RDATA_194;
   assign RDATA[1567:1560] = RDATA_195;
   assign RDATA[1575:1568] = RDATA_196;
   assign RDATA[1583:1576] = RDATA_197;
   assign RDATA[1591:1584] = RDATA_198;
   assign RDATA[1599:1592] = RDATA_199;
   assign RDATA[1607:1600] = RDATA_200;
   assign RDATA[1615:1608] = RDATA_201;
   assign RDATA[1623:1616] = RDATA_202;
   assign RDATA[1631:1624] = RDATA_203;
   assign RDATA[1639:1632] = RDATA_204;
   assign RDATA[1647:1640] = RDATA_205;
   assign RDATA[1655:1648] = RDATA_206;
   assign RDATA[1663:1656] = RDATA_207;
   assign RDATA[1671:1664] = RDATA_208;
   assign RDATA[1679:1672] = RDATA_209;
   assign RDATA[1687:1680] = RDATA_210;
   assign RDATA[1695:1688] = RDATA_211;
   assign RDATA[1703:1696] = RDATA_212;
   assign RDATA[1711:1704] = RDATA_213;
   assign RDATA[1719:1712] = RDATA_214;
   assign RDATA[1727:1720] = RDATA_215;
   assign RDATA[1735:1728] = RDATA_216;
   assign RDATA[1743:1736] = RDATA_217;
   assign RDATA[1751:1744] = RDATA_218;
   assign RDATA[1759:1752] = RDATA_219;
   assign RDATA[1767:1760] = RDATA_220;
   assign RDATA[1775:1768] = RDATA_221;
   assign RDATA[1783:1776] = RDATA_222;
   assign RDATA[1791:1784] = RDATA_223;
   assign RDATA[1799:1792] = RDATA_224;
   assign RDATA[1807:1800] = RDATA_225;
   assign RDATA[1815:1808] = RDATA_226;
   assign RDATA[1823:1816] = RDATA_227;
   assign RDATA[1831:1824] = RDATA_228;
   assign RDATA[1839:1832] = RDATA_229;
   assign RDATA[1847:1840] = RDATA_230;
   assign RDATA[1855:1848] = RDATA_231;
   assign RDATA[1863:1856] = RDATA_232;
   assign RDATA[1871:1864] = RDATA_233;
   assign RDATA[1879:1872] = RDATA_234;
   assign RDATA[1887:1880] = RDATA_235;
   assign RDATA[1895:1888] = RDATA_236;
   assign RDATA[1903:1896] = RDATA_237;
   assign RDATA[1911:1904] = RDATA_238;
   assign RDATA[1919:1912] = RDATA_239;
   assign RDATA[1927:1920] = RDATA_240;
   assign RDATA[1935:1928] = RDATA_241;
   assign RDATA[1943:1936] = RDATA_242;
   assign RDATA[1951:1944] = RDATA_243;
   assign RDATA[1959:1952] = RDATA_244;
   assign RDATA[1967:1960] = RDATA_245;
   assign RDATA[1975:1968] = RDATA_246;
   assign RDATA[1983:1976] = RDATA_247;
   assign RDATA[1991:1984] = RDATA_248;
   assign RDATA[1999:1992] = RDATA_249;
   assign RDATA[2007:2000] = RDATA_250;
   assign RDATA[2015:2008] = RDATA_251;
   assign RDATA[2023:2016] = RDATA_252;
   assign RDATA[2031:2024] = RDATA_253;
   assign RDATA[2039:2032] = RDATA_254;
   assign RDATA[2047:2040] = RDATA_255;
   assign RDATA[2055:2048] = RDATA_256;
   assign RDATA[2063:2056] = RDATA_257;
   assign RDATA[2071:2064] = RDATA_258;
   assign RDATA[2079:2072] = RDATA_259;
   assign RDATA[2087:2080] = RDATA_260;
   assign RDATA[2095:2088] = RDATA_261;
   assign RDATA[2103:2096] = RDATA_262;
   assign RDATA[2111:2104] = RDATA_263;
   assign RDATA[2119:2112] = RDATA_264;
   assign RDATA[2127:2120] = RDATA_265;
   assign RDATA[2135:2128] = RDATA_266;
   assign RDATA[2143:2136] = RDATA_267;
   assign RDATA[2151:2144] = RDATA_268;
   assign RDATA[2159:2152] = RDATA_269;
   assign RDATA[2167:2160] = RDATA_270;
   assign RDATA[2175:2168] = RDATA_271;
   assign RDATA[2183:2176] = RDATA_272;
   assign RDATA[2191:2184] = RDATA_273;
   assign RDATA[2199:2192] = RDATA_274;
   assign RDATA[2207:2200] = RDATA_275;
   assign RDATA[2215:2208] = RDATA_276;
   assign RDATA[2223:2216] = RDATA_277;
   assign RDATA[2231:2224] = RDATA_278;
   assign RDATA[2239:2232] = RDATA_279;
   assign RDATA[2247:2240] = RDATA_280;
   assign RDATA[2255:2248] = RDATA_281;
   assign RDATA[2263:2256] = RDATA_282;
   assign RDATA[2271:2264] = RDATA_283;
   assign RDATA[2279:2272] = RDATA_284;
   assign RDATA[2287:2280] = RDATA_285;
   assign RDATA[2295:2288] = RDATA_286;
   assign RDATA[2303:2296] = RDATA_287;
   assign RDATA[2311:2304] = RDATA_288;
   assign RDATA[2319:2312] = RDATA_289;
   assign RDATA[2327:2320] = RDATA_290;
   assign RDATA[2335:2328] = RDATA_291;
   assign RDATA[2343:2336] = RDATA_292;
   assign RDATA[2351:2344] = RDATA_293;
   assign RDATA[2359:2352] = RDATA_294;
   assign RDATA[2367:2360] = RDATA_295;
   assign RDATA[2375:2368] = RDATA_296;
   assign RDATA[2383:2376] = RDATA_297;
   assign RDATA[2391:2384] = RDATA_298;
   assign RDATA[2399:2392] = RDATA_299;
   assign RDATA[2407:2400] = RDATA_300;
   assign RDATA[2415:2408] = RDATA_301;
   assign RDATA[2423:2416] = RDATA_302;
   assign RDATA[2431:2424] = RDATA_303;
   assign RDATA[2439:2432] = RDATA_304;
   assign RDATA[2447:2440] = RDATA_305;
   assign RDATA[2455:2448] = RDATA_306;
   assign RDATA[2463:2456] = RDATA_307;
   assign RDATA[2471:2464] = RDATA_308;
   assign RDATA[2479:2472] = RDATA_309;
   assign RDATA[2487:2480] = RDATA_310;
   assign RDATA[2495:2488] = RDATA_311;
   assign RDATA[2503:2496] = RDATA_312;
   assign RDATA[2511:2504] = RDATA_313;
   assign RDATA[2519:2512] = RDATA_314;
   assign RDATA[2527:2520] = RDATA_315;
   assign RDATA[2535:2528] = RDATA_316;
   assign RDATA[2543:2536] = RDATA_317;
   assign RDATA[2551:2544] = RDATA_318;
   assign RDATA[2559:2552] = RDATA_319;
   assign RDATA[2567:2560] = RDATA_320;
   assign RDATA[2575:2568] = RDATA_321;
   assign RDATA[2583:2576] = RDATA_322;
   assign RDATA[2591:2584] = RDATA_323;
   assign RDATA[2599:2592] = RDATA_324;
   assign RDATA[2607:2600] = RDATA_325;
   assign RDATA[2615:2608] = RDATA_326;
   assign RDATA[2623:2616] = RDATA_327;
   assign RDATA[2631:2624] = RDATA_328;
   assign RDATA[2639:2632] = RDATA_329;
   assign RDATA[2647:2640] = RDATA_330;
   assign RDATA[2655:2648] = RDATA_331;
   assign RDATA[2663:2656] = RDATA_332;
   assign RDATA[2671:2664] = RDATA_333;
   assign RDATA[2679:2672] = RDATA_334;
   assign RDATA[2687:2680] = RDATA_335;
   assign RDATA[2695:2688] = RDATA_336;
   assign RDATA[2703:2696] = RDATA_337;
   assign RDATA[2711:2704] = RDATA_338;
   assign RDATA[2719:2712] = RDATA_339;
   assign RDATA[2727:2720] = RDATA_340;
   assign RDATA[2735:2728] = RDATA_341;
   assign RDATA[2743:2736] = RDATA_342;
   assign RDATA[2751:2744] = RDATA_343;
   assign RDATA[2759:2752] = RDATA_344;
   assign RDATA[2767:2760] = RDATA_345;
   assign RDATA[2775:2768] = RDATA_346;
   assign RDATA[2783:2776] = RDATA_347;
   assign RDATA[2791:2784] = RDATA_348;
   assign RDATA[2799:2792] = RDATA_349;
   assign RDATA[2807:2800] = RDATA_350;
   assign RDATA[2815:2808] = RDATA_351;
   assign RDATA[2823:2816] = RDATA_352;
   assign RDATA[2831:2824] = RDATA_353;
   assign RDATA[2839:2832] = RDATA_354;
   assign RDATA[2847:2840] = RDATA_355;
   assign RDATA[2855:2848] = RDATA_356;
   assign RDATA[2863:2856] = RDATA_357;
   assign RDATA[2871:2864] = RDATA_358;
   assign RDATA[2879:2872] = RDATA_359;
   assign RDATA[2887:2880] = RDATA_360;
   assign RDATA[2895:2888] = RDATA_361;
   assign RDATA[2903:2896] = RDATA_362;
   assign RDATA[2911:2904] = RDATA_363;
   assign RDATA[2919:2912] = RDATA_364;
   assign RDATA[2927:2920] = RDATA_365;
   assign RDATA[2935:2928] = RDATA_366;
   assign RDATA[2943:2936] = RDATA_367;
   assign RDATA[2951:2944] = RDATA_368;
   assign RDATA[2959:2952] = RDATA_369;
   assign RDATA[2967:2960] = RDATA_370;
   assign RDATA[2975:2968] = RDATA_371;
   assign RDATA[2983:2976] = RDATA_372;
   assign RDATA[2991:2984] = RDATA_373;
   assign RDATA[2999:2992] = RDATA_374;
   assign RDATA[3007:3000] = RDATA_375;
   assign RDATA[3015:3008] = RDATA_376;
   assign RDATA[3023:3016] = RDATA_377;
   assign RDATA[3031:3024] = RDATA_378;
   assign RDATA[3039:3032] = RDATA_379;
   assign RDATA[3047:3040] = RDATA_380;
   assign RDATA[3055:3048] = RDATA_381;
   assign RDATA[3063:3056] = RDATA_382;
   assign RDATA[3071:3064] = RDATA_383;
   assign RDATA[3079:3072] = RDATA_384;
   assign RDATA[3087:3080] = RDATA_385;
   assign RDATA[3095:3088] = RDATA_386;
   assign RDATA[3103:3096] = RDATA_387;
   assign RDATA[3111:3104] = RDATA_388;
   assign RDATA[3119:3112] = RDATA_389;
   assign RDATA[3127:3120] = RDATA_390;
   assign RDATA[3135:3128] = RDATA_391;
   assign RDATA[3143:3136] = RDATA_392;
   assign RDATA[3151:3144] = RDATA_393;
   assign RDATA[3159:3152] = RDATA_394;
   assign RDATA[3167:3160] = RDATA_395;
   assign RDATA[3175:3168] = RDATA_396;
   assign RDATA[3183:3176] = RDATA_397;
   assign RDATA[3191:3184] = RDATA_398;
   assign RDATA[3199:3192] = RDATA_399;
   assign RDATA[3207:3200] = RDATA_400;
   assign RDATA[3215:3208] = RDATA_401;
   assign RDATA[3223:3216] = RDATA_402;
   assign RDATA[3231:3224] = RDATA_403;
   assign RDATA[3239:3232] = RDATA_404;
   assign RDATA[3247:3240] = RDATA_405;
   assign RDATA[3255:3248] = RDATA_406;
   assign RDATA[3263:3256] = RDATA_407;
   assign RDATA[3271:3264] = RDATA_408;
   assign RDATA[3279:3272] = RDATA_409;
   assign RDATA[3287:3280] = RDATA_410;
   assign RDATA[3295:3288] = RDATA_411;
   assign RDATA[3303:3296] = RDATA_412;
   assign RDATA[3311:3304] = RDATA_413;
   assign RDATA[3319:3312] = RDATA_414;
   assign RDATA[3327:3320] = RDATA_415;
   assign RDATA[3335:3328] = RDATA_416;
   assign RDATA[3343:3336] = RDATA_417;
   assign RDATA[3351:3344] = RDATA_418;
   assign RDATA[3359:3352] = RDATA_419;
   assign RDATA[3367:3360] = RDATA_420;
   assign RDATA[3375:3368] = RDATA_421;
   assign RDATA[3383:3376] = RDATA_422;
   assign RDATA[3391:3384] = RDATA_423;
   assign RDATA[3399:3392] = RDATA_424;
   assign RDATA[3407:3400] = RDATA_425;
   assign RDATA[3415:3408] = RDATA_426;
   assign RDATA[3423:3416] = RDATA_427;
   assign RDATA[3431:3424] = RDATA_428;
   assign RDATA[3439:3432] = RDATA_429;
   assign RDATA[3447:3440] = RDATA_430;
   assign RDATA[3455:3448] = RDATA_431;
   assign RDATA[3463:3456] = RDATA_432;
   assign RDATA[3471:3464] = RDATA_433;
   assign RDATA[3479:3472] = RDATA_434;
   assign RDATA[3487:3480] = RDATA_435;
   assign RDATA[3495:3488] = RDATA_436;
   assign RDATA[3503:3496] = RDATA_437;
   assign RDATA[3511:3504] = RDATA_438;
   assign RDATA[3519:3512] = RDATA_439;
   assign RDATA[3527:3520] = RDATA_440;
   assign RDATA[3535:3528] = RDATA_441;
   assign RDATA[3543:3536] = RDATA_442;
   assign RDATA[3551:3544] = RDATA_443;
   assign RDATA[3559:3552] = RDATA_444;
   assign RDATA[3567:3560] = RDATA_445;
   assign RDATA[3575:3568] = RDATA_446;
   assign RDATA[3583:3576] = RDATA_447;
   assign RDATA[3591:3584] = RDATA_448;
   assign RDATA[3599:3592] = RDATA_449;
   assign RDATA[3607:3600] = RDATA_450;
   assign RDATA[3615:3608] = RDATA_451;
   assign RDATA[3623:3616] = RDATA_452;
   assign RDATA[3631:3624] = RDATA_453;
   assign RDATA[3639:3632] = RDATA_454;
   assign RDATA[3647:3640] = RDATA_455;
   assign RDATA[3655:3648] = RDATA_456;
   assign RDATA[3663:3656] = RDATA_457;
   assign RDATA[3671:3664] = RDATA_458;
   assign RDATA[3679:3672] = RDATA_459;
   assign RDATA[3687:3680] = RDATA_460;
   assign RDATA[3695:3688] = RDATA_461;
   assign RDATA[3703:3696] = RDATA_462;
   assign RDATA[3711:3704] = RDATA_463;
   assign RDATA[3719:3712] = RDATA_464;
   assign RDATA[3727:3720] = RDATA_465;
   assign RDATA[3735:3728] = RDATA_466;
   assign RDATA[3743:3736] = RDATA_467;
   assign RDATA[3751:3744] = RDATA_468;
   assign RDATA[3759:3752] = RDATA_469;
   assign RDATA[3767:3760] = RDATA_470;
   assign RDATA[3775:3768] = RDATA_471;
   assign RDATA[3783:3776] = RDATA_472;
   assign RDATA[3791:3784] = RDATA_473;
   assign RDATA[3799:3792] = RDATA_474;
   assign RDATA[3807:3800] = RDATA_475;
   assign RDATA[3815:3808] = RDATA_476;
   assign RDATA[3823:3816] = RDATA_477;
   assign RDATA[3831:3824] = RDATA_478;
   assign RDATA[3839:3832] = RDATA_479;
   assign RDATA[3847:3840] = RDATA_480;
   assign RDATA[3855:3848] = RDATA_481;
   assign RDATA[3863:3856] = RDATA_482;
   assign RDATA[3871:3864] = RDATA_483;
   assign RDATA[3879:3872] = RDATA_484;
   assign RDATA[3887:3880] = RDATA_485;
   assign RDATA[3895:3888] = RDATA_486;
   assign RDATA[3903:3896] = RDATA_487;
   assign RDATA[3911:3904] = RDATA_488;
   assign RDATA[3919:3912] = RDATA_489;
   assign RDATA[3927:3920] = RDATA_490;
   assign RDATA[3935:3928] = RDATA_491;
   assign RDATA[3943:3936] = RDATA_492;
   assign RDATA[3951:3944] = RDATA_493;
   assign RDATA[3959:3952] = RDATA_494;
   assign RDATA[3967:3960] = RDATA_495;
   assign RDATA[3975:3968] = RDATA_496;
   assign RDATA[3983:3976] = RDATA_497;
   assign RDATA[3991:3984] = RDATA_498;
   assign RDATA[3999:3992] = RDATA_499;
   assign RDATA[4007:4000] = RDATA_500;
   assign RDATA[4015:4008] = RDATA_501;
   assign RDATA[4023:4016] = RDATA_502;
   assign RDATA[4031:4024] = RDATA_503;
   assign RDATA[4039:4032] = RDATA_504;
   assign RDATA[4047:4040] = RDATA_505;
   assign RDATA[4055:4048] = RDATA_506;
   assign RDATA[4063:4056] = RDATA_507;
   assign RDATA[4071:4064] = RDATA_508;
   assign RDATA[4079:4072] = RDATA_509;
   assign RDATA[4087:4080] = RDATA_510;
   assign RDATA[4095:4088] = RDATA_511;
   assign RDATA[4103:4096] = RDATA_512;
   assign RDATA[4111:4104] = RDATA_513;
   assign RDATA[4119:4112] = RDATA_514;
   assign RDATA[4127:4120] = RDATA_515;
   assign RDATA[4135:4128] = RDATA_516;
   assign RDATA[4143:4136] = RDATA_517;
   assign RDATA[4151:4144] = RDATA_518;
   assign RDATA[4159:4152] = RDATA_519;
   assign RDATA[4167:4160] = RDATA_520;
   assign RDATA[4175:4168] = RDATA_521;
   assign RDATA[4183:4176] = RDATA_522;
   assign RDATA[4191:4184] = RDATA_523;
   assign RDATA[4199:4192] = RDATA_524;
   assign RDATA[4207:4200] = RDATA_525;
   assign RDATA[4215:4208] = RDATA_526;
   assign RDATA[4223:4216] = RDATA_527;
   assign RDATA[4231:4224] = RDATA_528;
   assign RDATA[4239:4232] = RDATA_529;
   assign RDATA[4247:4240] = RDATA_530;
   assign RDATA[4255:4248] = RDATA_531;
   assign RDATA[4263:4256] = RDATA_532;
   assign RDATA[4271:4264] = RDATA_533;
   assign RDATA[4279:4272] = RDATA_534;
   assign RDATA[4287:4280] = RDATA_535;
   assign RDATA[4295:4288] = RDATA_536;
   assign RDATA[4303:4296] = RDATA_537;
   assign RDATA[4311:4304] = RDATA_538;
   assign RDATA[4319:4312] = RDATA_539;
   assign RDATA[4327:4320] = RDATA_540;
   assign RDATA[4335:4328] = RDATA_541;
   assign RDATA[4343:4336] = RDATA_542;
   assign RDATA[4351:4344] = RDATA_543;
   assign RDATA[4359:4352] = RDATA_544;
   assign RDATA[4367:4360] = RDATA_545;
   assign RDATA[4375:4368] = RDATA_546;
   assign RDATA[4383:4376] = RDATA_547;
   assign RDATA[4391:4384] = RDATA_548;
   assign RDATA[4399:4392] = RDATA_549;
   assign RDATA[4407:4400] = RDATA_550;
   assign RDATA[4415:4408] = RDATA_551;
   assign RDATA[4423:4416] = RDATA_552;
   assign RDATA[4431:4424] = RDATA_553;
   assign RDATA[4439:4432] = RDATA_554;
   assign RDATA[4447:4440] = RDATA_555;
   assign RDATA[4455:4448] = RDATA_556;
   assign RDATA[4463:4456] = RDATA_557;
   assign RDATA[4471:4464] = RDATA_558;
   assign RDATA[4479:4472] = RDATA_559;
   assign RDATA[4487:4480] = RDATA_560;
   assign RDATA[4495:4488] = RDATA_561;
   assign RDATA[4503:4496] = RDATA_562;
   assign RDATA[4511:4504] = RDATA_563;
   assign RDATA[4519:4512] = RDATA_564;
   assign RDATA[4527:4520] = RDATA_565;
   assign RDATA[4535:4528] = RDATA_566;
   assign RDATA[4543:4536] = RDATA_567;
   assign RDATA[4551:4544] = RDATA_568;
   assign RDATA[4559:4552] = RDATA_569;
   assign RDATA[4567:4560] = RDATA_570;
   assign RDATA[4575:4568] = RDATA_571;
   assign RDATA[4583:4576] = RDATA_572;
   assign RDATA[4591:4584] = RDATA_573;
   assign RDATA[4599:4592] = RDATA_574;
   assign RDATA[4607:4600] = RDATA_575;
   assign RDATA[4615:4608] = RDATA_576;
   assign RDATA[4623:4616] = RDATA_577;
   assign RDATA[4631:4624] = RDATA_578;
   assign RDATA[4639:4632] = RDATA_579;
   assign RDATA[4647:4640] = RDATA_580;
   assign RDATA[4655:4648] = RDATA_581;
   assign RDATA[4663:4656] = RDATA_582;
   assign RDATA[4671:4664] = RDATA_583;
   assign RDATA[4679:4672] = RDATA_584;
   assign RDATA[4687:4680] = RDATA_585;
   assign RDATA[4695:4688] = RDATA_586;
   assign RDATA[4703:4696] = RDATA_587;
   assign RDATA[4711:4704] = RDATA_588;
   assign RDATA[4719:4712] = RDATA_589;
   assign RDATA[4727:4720] = RDATA_590;
   assign RDATA[4735:4728] = RDATA_591;
   assign RDATA[4743:4736] = RDATA_592;
   assign RDATA[4751:4744] = RDATA_593;
   assign RDATA[4759:4752] = RDATA_594;
   assign RDATA[4767:4760] = RDATA_595;
   assign RDATA[4775:4768] = RDATA_596;
   assign RDATA[4783:4776] = RDATA_597;
   assign RDATA[4791:4784] = RDATA_598;
   assign RDATA[4799:4792] = RDATA_599;
   assign RDATA[4807:4800] = RDATA_600;
   assign RDATA[4815:4808] = RDATA_601;
   assign RDATA[4823:4816] = RDATA_602;
   assign RDATA[4831:4824] = RDATA_603;
   assign RDATA[4839:4832] = RDATA_604;
   assign RDATA[4847:4840] = RDATA_605;
   assign RDATA[4855:4848] = RDATA_606;
   assign RDATA[4863:4856] = RDATA_607;
   assign RDATA[4871:4864] = RDATA_608;
   assign RDATA[4879:4872] = RDATA_609;
   assign RDATA[4887:4880] = RDATA_610;
   assign RDATA[4895:4888] = RDATA_611;
   assign RDATA[4903:4896] = RDATA_612;
   assign RDATA[4911:4904] = RDATA_613;
   assign RDATA[4919:4912] = RDATA_614;
   assign RDATA[4927:4920] = RDATA_615;
   assign RDATA[4935:4928] = RDATA_616;
   assign RDATA[4943:4936] = RDATA_617;
   assign RDATA[4951:4944] = RDATA_618;
   assign RDATA[4959:4952] = RDATA_619;
   assign RDATA[4967:4960] = RDATA_620;
   assign RDATA[4975:4968] = RDATA_621;
   assign RDATA[4983:4976] = RDATA_622;
   assign RDATA[4991:4984] = RDATA_623;
   assign RDATA[4999:4992] = RDATA_624;
   assign RDATA[5007:5000] = RDATA_625;
   assign RDATA[5015:5008] = RDATA_626;
   assign RDATA[5023:5016] = RDATA_627;
   assign RDATA[5031:5024] = RDATA_628;
   assign RDATA[5039:5032] = RDATA_629;
   assign RDATA[5047:5040] = RDATA_630;
   assign RDATA[5055:5048] = RDATA_631;
   assign RDATA[5063:5056] = RDATA_632;
   assign RDATA[5071:5064] = RDATA_633;
   assign RDATA[5079:5072] = RDATA_634;
   assign RDATA[5087:5080] = RDATA_635;
   assign RDATA[5095:5088] = RDATA_636;
   assign RDATA[5103:5096] = RDATA_637;
   assign RDATA[5111:5104] = RDATA_638;
   assign RDATA[5119:5112] = RDATA_639;
   assign RDATA[5127:5120] = RDATA_640;
   assign RDATA[5135:5128] = RDATA_641;
   assign RDATA[5143:5136] = RDATA_642;
   assign RDATA[5151:5144] = RDATA_643;
   assign RDATA[5159:5152] = RDATA_644;
   assign RDATA[5167:5160] = RDATA_645;
   assign RDATA[5175:5168] = RDATA_646;
   assign RDATA[5183:5176] = RDATA_647;
   assign RDATA[5191:5184] = RDATA_648;
   assign RDATA[5199:5192] = RDATA_649;
   assign RDATA[5207:5200] = RDATA_650;
   assign RDATA[5215:5208] = RDATA_651;
   assign RDATA[5223:5216] = RDATA_652;
   assign RDATA[5231:5224] = RDATA_653;
   assign RDATA[5239:5232] = RDATA_654;
   assign RDATA[5247:5240] = RDATA_655;
   assign RDATA[5255:5248] = RDATA_656;
   assign RDATA[5263:5256] = RDATA_657;
   assign RDATA[5271:5264] = RDATA_658;
   assign RDATA[5279:5272] = RDATA_659;
   assign RDATA[5287:5280] = RDATA_660;
   assign RDATA[5295:5288] = RDATA_661;
   assign RDATA[5303:5296] = RDATA_662;
   assign RDATA[5311:5304] = RDATA_663;
   assign RDATA[5319:5312] = RDATA_664;
   assign RDATA[5327:5320] = RDATA_665;
   assign RDATA[5335:5328] = RDATA_666;
   assign RDATA[5343:5336] = RDATA_667;
   assign RDATA[5351:5344] = RDATA_668;
   assign RDATA[5359:5352] = RDATA_669;
   assign RDATA[5367:5360] = RDATA_670;
   assign RDATA[5375:5368] = RDATA_671;
   assign RDATA[5383:5376] = RDATA_672;
   assign RDATA[5391:5384] = RDATA_673;
   assign RDATA[5399:5392] = RDATA_674;
   assign RDATA[5407:5400] = RDATA_675;
   assign RDATA[5415:5408] = RDATA_676;
   assign RDATA[5423:5416] = RDATA_677;
   assign RDATA[5431:5424] = RDATA_678;
   assign RDATA[5439:5432] = RDATA_679;
   assign RDATA[5447:5440] = RDATA_680;
   assign RDATA[5455:5448] = RDATA_681;
   assign RDATA[5463:5456] = RDATA_682;
   assign RDATA[5471:5464] = RDATA_683;
   assign RDATA[5479:5472] = RDATA_684;
   assign RDATA[5487:5480] = RDATA_685;
   assign RDATA[5495:5488] = RDATA_686;
   assign RDATA[5503:5496] = RDATA_687;
   assign RDATA[5511:5504] = RDATA_688;
   assign RDATA[5519:5512] = RDATA_689;
   assign RDATA[5527:5520] = RDATA_690;
   assign RDATA[5535:5528] = RDATA_691;
   assign RDATA[5543:5536] = RDATA_692;
   assign RDATA[5551:5544] = RDATA_693;
   assign RDATA[5559:5552] = RDATA_694;
   assign RDATA[5567:5560] = RDATA_695;
   assign RDATA[5575:5568] = RDATA_696;
   assign RDATA[5583:5576] = RDATA_697;
   assign RDATA[5591:5584] = RDATA_698;
   assign RDATA[5599:5592] = RDATA_699;
   assign RDATA[5607:5600] = RDATA_700;
   assign RDATA[5615:5608] = RDATA_701;
   assign RDATA[5623:5616] = RDATA_702;
   assign RDATA[5631:5624] = RDATA_703;
   assign RDATA[5639:5632] = RDATA_704;
   assign RDATA[5647:5640] = RDATA_705;
   assign RDATA[5655:5648] = RDATA_706;
   assign RDATA[5663:5656] = RDATA_707;
   assign RDATA[5671:5664] = RDATA_708;
   assign RDATA[5679:5672] = RDATA_709;
   assign RDATA[5687:5680] = RDATA_710;
   assign RDATA[5695:5688] = RDATA_711;
   assign RDATA[5703:5696] = RDATA_712;
   assign RDATA[5711:5704] = RDATA_713;
   assign RDATA[5719:5712] = RDATA_714;
   assign RDATA[5727:5720] = RDATA_715;
   assign RDATA[5735:5728] = RDATA_716;
   assign RDATA[5743:5736] = RDATA_717;
   assign RDATA[5751:5744] = RDATA_718;
   assign RDATA[5759:5752] = RDATA_719;
   assign RDATA[5767:5760] = RDATA_720;
   assign RDATA[5775:5768] = RDATA_721;
   assign RDATA[5783:5776] = RDATA_722;
   assign RDATA[5791:5784] = RDATA_723;
   assign RDATA[5799:5792] = RDATA_724;
   assign RDATA[5807:5800] = RDATA_725;
   assign RDATA[5815:5808] = RDATA_726;
   assign RDATA[5823:5816] = RDATA_727;
   assign RDATA[5831:5824] = RDATA_728;
   assign RDATA[5839:5832] = RDATA_729;
   assign RDATA[5847:5840] = RDATA_730;
   assign RDATA[5855:5848] = RDATA_731;
   assign RDATA[5863:5856] = RDATA_732;
   assign RDATA[5871:5864] = RDATA_733;
   assign RDATA[5879:5872] = RDATA_734;
   assign RDATA[5887:5880] = RDATA_735;
   assign RDATA[5895:5888] = RDATA_736;
   assign RDATA[5903:5896] = RDATA_737;
   assign RDATA[5911:5904] = RDATA_738;
   assign RDATA[5919:5912] = RDATA_739;
   assign RDATA[5927:5920] = RDATA_740;
   assign RDATA[5935:5928] = RDATA_741;
   assign RDATA[5943:5936] = RDATA_742;
   assign RDATA[5951:5944] = RDATA_743;
   assign RDATA[5959:5952] = RDATA_744;
   assign RDATA[5967:5960] = RDATA_745;
   assign RDATA[5975:5968] = RDATA_746;
   assign RDATA[5983:5976] = RDATA_747;
   assign RDATA[5991:5984] = RDATA_748;
   assign RDATA[5999:5992] = RDATA_749;
   assign RDATA[6007:6000] = RDATA_750;
   assign RDATA[6015:6008] = RDATA_751;
   assign RDATA[6023:6016] = RDATA_752;
   assign RDATA[6031:6024] = RDATA_753;
   assign RDATA[6039:6032] = RDATA_754;
   assign RDATA[6047:6040] = RDATA_755;
   assign RDATA[6055:6048] = RDATA_756;
   assign RDATA[6063:6056] = RDATA_757;
   assign RDATA[6071:6064] = RDATA_758;
   assign RDATA[6079:6072] = RDATA_759;
   assign RDATA[6087:6080] = RDATA_760;
   assign RDATA[6095:6088] = RDATA_761;
   assign RDATA[6103:6096] = RDATA_762;
   assign RDATA[6111:6104] = RDATA_763;
   assign RDATA[6119:6112] = RDATA_764;
   assign RDATA[6127:6120] = RDATA_765;
   assign RDATA[6135:6128] = RDATA_766;
   assign RDATA[6143:6136] = RDATA_767;
   assign RDATA[6151:6144] = RDATA_768;
   assign RDATA[6159:6152] = RDATA_769;
   assign RDATA[6167:6160] = RDATA_770;
   assign RDATA[6175:6168] = RDATA_771;
   assign RDATA[6183:6176] = RDATA_772;
   assign RDATA[6191:6184] = RDATA_773;
   assign RDATA[6199:6192] = RDATA_774;
   assign RDATA[6207:6200] = RDATA_775;
   assign RDATA[6215:6208] = RDATA_776;
   assign RDATA[6223:6216] = RDATA_777;
   assign RDATA[6231:6224] = RDATA_778;
   assign RDATA[6239:6232] = RDATA_779;
   assign RDATA[6247:6240] = RDATA_780;
   assign RDATA[6255:6248] = RDATA_781;
   assign RDATA[6263:6256] = RDATA_782;
   assign RDATA[6271:6264] = RDATA_783;

   

endmodule // img_sram
