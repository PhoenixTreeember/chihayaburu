module mul_add_core
  (
   input 	       CLK,
   input 	       RESET_X,

   input [28*28*8-1:0] W,
   input [7:0] 	       B,
   input [28*28*8-1:0] IMG,

   output reg [31:0]       RESULT
   
   );


   wire [7:0] 	       mul_out_0;
   wire [7:0] 	       mul_out_1;
   wire [7:0] 	       mul_out_2;
   wire [7:0] 	       mul_out_3;
   wire [7:0] 	       mul_out_4;
   wire [7:0] 	       mul_out_5;
   wire [7:0] 	       mul_out_6;
   wire [7:0] 	       mul_out_7;
   wire [7:0] 	       mul_out_8;
   wire [7:0] 	       mul_out_9;
   wire [7:0] 	       mul_out_10;
   wire [7:0] 	       mul_out_11;
   wire [7:0] 	       mul_out_12;
   wire [7:0] 	       mul_out_13;
   wire [7:0] 	       mul_out_14;
   wire [7:0] 	       mul_out_15;
   wire [7:0] 	       mul_out_16;
   wire [7:0] 	       mul_out_17;
   wire [7:0] 	       mul_out_18;
   wire [7:0] 	       mul_out_19;
   wire [7:0] 	       mul_out_20;
   wire [7:0] 	       mul_out_21;
   wire [7:0] 	       mul_out_22;
   wire [7:0] 	       mul_out_23;
   wire [7:0] 	       mul_out_24;
   wire [7:0] 	       mul_out_25;
   wire [7:0] 	       mul_out_26;
   wire [7:0] 	       mul_out_27;
   wire [7:0] 	       mul_out_28;
   wire [7:0] 	       mul_out_29;
   wire [7:0] 	       mul_out_30;
   wire [7:0] 	       mul_out_31;
   wire [7:0] 	       mul_out_32;
   wire [7:0] 	       mul_out_33;
   wire [7:0] 	       mul_out_34;
   wire [7:0] 	       mul_out_35;
   wire [7:0] 	       mul_out_36;
   wire [7:0] 	       mul_out_37;
   wire [7:0] 	       mul_out_38;
   wire [7:0] 	       mul_out_39;
   wire [7:0] 	       mul_out_40;
   wire [7:0] 	       mul_out_41;
   wire [7:0] 	       mul_out_42;
   wire [7:0] 	       mul_out_43;
   wire [7:0] 	       mul_out_44;
   wire [7:0] 	       mul_out_45;
   wire [7:0] 	       mul_out_46;
   wire [7:0] 	       mul_out_47;
   wire [7:0] 	       mul_out_48;
   wire [7:0] 	       mul_out_49;
   wire [7:0] 	       mul_out_50;
   wire [7:0] 	       mul_out_51;
   wire [7:0] 	       mul_out_52;
   wire [7:0] 	       mul_out_53;
   wire [7:0] 	       mul_out_54;
   wire [7:0] 	       mul_out_55;
   wire [7:0] 	       mul_out_56;
   wire [7:0] 	       mul_out_57;
   wire [7:0] 	       mul_out_58;
   wire [7:0] 	       mul_out_59;
   wire [7:0] 	       mul_out_60;
   wire [7:0] 	       mul_out_61;
   wire [7:0] 	       mul_out_62;
   wire [7:0] 	       mul_out_63;
   wire [7:0] 	       mul_out_64;
   wire [7:0] 	       mul_out_65;
   wire [7:0] 	       mul_out_66;
   wire [7:0] 	       mul_out_67;
   wire [7:0] 	       mul_out_68;
   wire [7:0] 	       mul_out_69;
   wire [7:0] 	       mul_out_70;
   wire [7:0] 	       mul_out_71;
   wire [7:0] 	       mul_out_72;
   wire [7:0] 	       mul_out_73;
   wire [7:0] 	       mul_out_74;
   wire [7:0] 	       mul_out_75;
   wire [7:0] 	       mul_out_76;
   wire [7:0] 	       mul_out_77;
   wire [7:0] 	       mul_out_78;
   wire [7:0] 	       mul_out_79;
   wire [7:0] 	       mul_out_80;
   wire [7:0] 	       mul_out_81;
   wire [7:0] 	       mul_out_82;
   wire [7:0] 	       mul_out_83;
   wire [7:0] 	       mul_out_84;
   wire [7:0] 	       mul_out_85;
   wire [7:0] 	       mul_out_86;
   wire [7:0] 	       mul_out_87;
   wire [7:0] 	       mul_out_88;
   wire [7:0] 	       mul_out_89;
   wire [7:0] 	       mul_out_90;
   wire [7:0] 	       mul_out_91;
   wire [7:0] 	       mul_out_92;
   wire [7:0] 	       mul_out_93;
   wire [7:0] 	       mul_out_94;
   wire [7:0] 	       mul_out_95;
   wire [7:0] 	       mul_out_96;
   wire [7:0] 	       mul_out_97;
   wire [7:0] 	       mul_out_98;
   wire [7:0] 	       mul_out_99;
   wire [7:0] 	       mul_out_100;
   wire [7:0] 	       mul_out_101;
   wire [7:0] 	       mul_out_102;
   wire [7:0] 	       mul_out_103;
   wire [7:0] 	       mul_out_104;
   wire [7:0] 	       mul_out_105;
   wire [7:0] 	       mul_out_106;
   wire [7:0] 	       mul_out_107;
   wire [7:0] 	       mul_out_108;
   wire [7:0] 	       mul_out_109;
   wire [7:0] 	       mul_out_110;
   wire [7:0] 	       mul_out_111;
   wire [7:0] 	       mul_out_112;
   wire [7:0] 	       mul_out_113;
   wire [7:0] 	       mul_out_114;
   wire [7:0] 	       mul_out_115;
   wire [7:0] 	       mul_out_116;
   wire [7:0] 	       mul_out_117;
   wire [7:0] 	       mul_out_118;
   wire [7:0] 	       mul_out_119;
   wire [7:0] 	       mul_out_120;
   wire [7:0] 	       mul_out_121;
   wire [7:0] 	       mul_out_122;
   wire [7:0] 	       mul_out_123;
   wire [7:0] 	       mul_out_124;
   wire [7:0] 	       mul_out_125;
   wire [7:0] 	       mul_out_126;
   wire [7:0] 	       mul_out_127;
   wire [7:0] 	       mul_out_128;
   wire [7:0] 	       mul_out_129;
   wire [7:0] 	       mul_out_130;
   wire [7:0] 	       mul_out_131;
   wire [7:0] 	       mul_out_132;
   wire [7:0] 	       mul_out_133;
   wire [7:0] 	       mul_out_134;
   wire [7:0] 	       mul_out_135;
   wire [7:0] 	       mul_out_136;
   wire [7:0] 	       mul_out_137;
   wire [7:0] 	       mul_out_138;
   wire [7:0] 	       mul_out_139;
   wire [7:0] 	       mul_out_140;
   wire [7:0] 	       mul_out_141;
   wire [7:0] 	       mul_out_142;
   wire [7:0] 	       mul_out_143;
   wire [7:0] 	       mul_out_144;
   wire [7:0] 	       mul_out_145;
   wire [7:0] 	       mul_out_146;
   wire [7:0] 	       mul_out_147;
   wire [7:0] 	       mul_out_148;
   wire [7:0] 	       mul_out_149;
   wire [7:0] 	       mul_out_150;
   wire [7:0] 	       mul_out_151;
   wire [7:0] 	       mul_out_152;
   wire [7:0] 	       mul_out_153;
   wire [7:0] 	       mul_out_154;
   wire [7:0] 	       mul_out_155;
   wire [7:0] 	       mul_out_156;
   wire [7:0] 	       mul_out_157;
   wire [7:0] 	       mul_out_158;
   wire [7:0] 	       mul_out_159;
   wire [7:0] 	       mul_out_160;
   wire [7:0] 	       mul_out_161;
   wire [7:0] 	       mul_out_162;
   wire [7:0] 	       mul_out_163;
   wire [7:0] 	       mul_out_164;
   wire [7:0] 	       mul_out_165;
   wire [7:0] 	       mul_out_166;
   wire [7:0] 	       mul_out_167;
   wire [7:0] 	       mul_out_168;
   wire [7:0] 	       mul_out_169;
   wire [7:0] 	       mul_out_170;
   wire [7:0] 	       mul_out_171;
   wire [7:0] 	       mul_out_172;
   wire [7:0] 	       mul_out_173;
   wire [7:0] 	       mul_out_174;
   wire [7:0] 	       mul_out_175;
   wire [7:0] 	       mul_out_176;
   wire [7:0] 	       mul_out_177;
   wire [7:0] 	       mul_out_178;
   wire [7:0] 	       mul_out_179;
   wire [7:0] 	       mul_out_180;
   wire [7:0] 	       mul_out_181;
   wire [7:0] 	       mul_out_182;
   wire [7:0] 	       mul_out_183;
   wire [7:0] 	       mul_out_184;
   wire [7:0] 	       mul_out_185;
   wire [7:0] 	       mul_out_186;
   wire [7:0] 	       mul_out_187;
   wire [7:0] 	       mul_out_188;
   wire [7:0] 	       mul_out_189;
   wire [7:0] 	       mul_out_190;
   wire [7:0] 	       mul_out_191;
   wire [7:0] 	       mul_out_192;
   wire [7:0] 	       mul_out_193;
   wire [7:0] 	       mul_out_194;
   wire [7:0] 	       mul_out_195;
   wire [7:0] 	       mul_out_196;
   wire [7:0] 	       mul_out_197;
   wire [7:0] 	       mul_out_198;
   wire [7:0] 	       mul_out_199;
   wire [7:0] 	       mul_out_200;
   wire [7:0] 	       mul_out_201;
   wire [7:0] 	       mul_out_202;
   wire [7:0] 	       mul_out_203;
   wire [7:0] 	       mul_out_204;
   wire [7:0] 	       mul_out_205;
   wire [7:0] 	       mul_out_206;
   wire [7:0] 	       mul_out_207;
   wire [7:0] 	       mul_out_208;
   wire [7:0] 	       mul_out_209;
   wire [7:0] 	       mul_out_210;
   wire [7:0] 	       mul_out_211;
   wire [7:0] 	       mul_out_212;
   wire [7:0] 	       mul_out_213;
   wire [7:0] 	       mul_out_214;
   wire [7:0] 	       mul_out_215;
   wire [7:0] 	       mul_out_216;
   wire [7:0] 	       mul_out_217;
   wire [7:0] 	       mul_out_218;
   wire [7:0] 	       mul_out_219;
   wire [7:0] 	       mul_out_220;
   wire [7:0] 	       mul_out_221;
   wire [7:0] 	       mul_out_222;
   wire [7:0] 	       mul_out_223;
   wire [7:0] 	       mul_out_224;
   wire [7:0] 	       mul_out_225;
   wire [7:0] 	       mul_out_226;
   wire [7:0] 	       mul_out_227;
   wire [7:0] 	       mul_out_228;
   wire [7:0] 	       mul_out_229;
   wire [7:0] 	       mul_out_230;
   wire [7:0] 	       mul_out_231;
   wire [7:0] 	       mul_out_232;
   wire [7:0] 	       mul_out_233;
   wire [7:0] 	       mul_out_234;
   wire [7:0] 	       mul_out_235;
   wire [7:0] 	       mul_out_236;
   wire [7:0] 	       mul_out_237;
   wire [7:0] 	       mul_out_238;
   wire [7:0] 	       mul_out_239;
   wire [7:0] 	       mul_out_240;
   wire [7:0] 	       mul_out_241;
   wire [7:0] 	       mul_out_242;
   wire [7:0] 	       mul_out_243;
   wire [7:0] 	       mul_out_244;
   wire [7:0] 	       mul_out_245;
   wire [7:0] 	       mul_out_246;
   wire [7:0] 	       mul_out_247;
   wire [7:0] 	       mul_out_248;
   wire [7:0] 	       mul_out_249;
   wire [7:0] 	       mul_out_250;
   wire [7:0] 	       mul_out_251;
   wire [7:0] 	       mul_out_252;
   wire [7:0] 	       mul_out_253;
   wire [7:0] 	       mul_out_254;
   wire [7:0] 	       mul_out_255;
   wire [7:0] 	       mul_out_256;
   wire [7:0] 	       mul_out_257;
   wire [7:0] 	       mul_out_258;
   wire [7:0] 	       mul_out_259;
   wire [7:0] 	       mul_out_260;
   wire [7:0] 	       mul_out_261;
   wire [7:0] 	       mul_out_262;
   wire [7:0] 	       mul_out_263;
   wire [7:0] 	       mul_out_264;
   wire [7:0] 	       mul_out_265;
   wire [7:0] 	       mul_out_266;
   wire [7:0] 	       mul_out_267;
   wire [7:0] 	       mul_out_268;
   wire [7:0] 	       mul_out_269;
   wire [7:0] 	       mul_out_270;
   wire [7:0] 	       mul_out_271;
   wire [7:0] 	       mul_out_272;
   wire [7:0] 	       mul_out_273;
   wire [7:0] 	       mul_out_274;
   wire [7:0] 	       mul_out_275;
   wire [7:0] 	       mul_out_276;
   wire [7:0] 	       mul_out_277;
   wire [7:0] 	       mul_out_278;
   wire [7:0] 	       mul_out_279;
   wire [7:0] 	       mul_out_280;
   wire [7:0] 	       mul_out_281;
   wire [7:0] 	       mul_out_282;
   wire [7:0] 	       mul_out_283;
   wire [7:0] 	       mul_out_284;
   wire [7:0] 	       mul_out_285;
   wire [7:0] 	       mul_out_286;
   wire [7:0] 	       mul_out_287;
   wire [7:0] 	       mul_out_288;
   wire [7:0] 	       mul_out_289;
   wire [7:0] 	       mul_out_290;
   wire [7:0] 	       mul_out_291;
   wire [7:0] 	       mul_out_292;
   wire [7:0] 	       mul_out_293;
   wire [7:0] 	       mul_out_294;
   wire [7:0] 	       mul_out_295;
   wire [7:0] 	       mul_out_296;
   wire [7:0] 	       mul_out_297;
   wire [7:0] 	       mul_out_298;
   wire [7:0] 	       mul_out_299;
   wire [7:0] 	       mul_out_300;
   wire [7:0] 	       mul_out_301;
   wire [7:0] 	       mul_out_302;
   wire [7:0] 	       mul_out_303;
   wire [7:0] 	       mul_out_304;
   wire [7:0] 	       mul_out_305;
   wire [7:0] 	       mul_out_306;
   wire [7:0] 	       mul_out_307;
   wire [7:0] 	       mul_out_308;
   wire [7:0] 	       mul_out_309;
   wire [7:0] 	       mul_out_310;
   wire [7:0] 	       mul_out_311;
   wire [7:0] 	       mul_out_312;
   wire [7:0] 	       mul_out_313;
   wire [7:0] 	       mul_out_314;
   wire [7:0] 	       mul_out_315;
   wire [7:0] 	       mul_out_316;
   wire [7:0] 	       mul_out_317;
   wire [7:0] 	       mul_out_318;
   wire [7:0] 	       mul_out_319;
   wire [7:0] 	       mul_out_320;
   wire [7:0] 	       mul_out_321;
   wire [7:0] 	       mul_out_322;
   wire [7:0] 	       mul_out_323;
   wire [7:0] 	       mul_out_324;
   wire [7:0] 	       mul_out_325;
   wire [7:0] 	       mul_out_326;
   wire [7:0] 	       mul_out_327;
   wire [7:0] 	       mul_out_328;
   wire [7:0] 	       mul_out_329;
   wire [7:0] 	       mul_out_330;
   wire [7:0] 	       mul_out_331;
   wire [7:0] 	       mul_out_332;
   wire [7:0] 	       mul_out_333;
   wire [7:0] 	       mul_out_334;
   wire [7:0] 	       mul_out_335;
   wire [7:0] 	       mul_out_336;
   wire [7:0] 	       mul_out_337;
   wire [7:0] 	       mul_out_338;
   wire [7:0] 	       mul_out_339;
   wire [7:0] 	       mul_out_340;
   wire [7:0] 	       mul_out_341;
   wire [7:0] 	       mul_out_342;
   wire [7:0] 	       mul_out_343;
   wire [7:0] 	       mul_out_344;
   wire [7:0] 	       mul_out_345;
   wire [7:0] 	       mul_out_346;
   wire [7:0] 	       mul_out_347;
   wire [7:0] 	       mul_out_348;
   wire [7:0] 	       mul_out_349;
   wire [7:0] 	       mul_out_350;
   wire [7:0] 	       mul_out_351;
   wire [7:0] 	       mul_out_352;
   wire [7:0] 	       mul_out_353;
   wire [7:0] 	       mul_out_354;
   wire [7:0] 	       mul_out_355;
   wire [7:0] 	       mul_out_356;
   wire [7:0] 	       mul_out_357;
   wire [7:0] 	       mul_out_358;
   wire [7:0] 	       mul_out_359;
   wire [7:0] 	       mul_out_360;
   wire [7:0] 	       mul_out_361;
   wire [7:0] 	       mul_out_362;
   wire [7:0] 	       mul_out_363;
   wire [7:0] 	       mul_out_364;
   wire [7:0] 	       mul_out_365;
   wire [7:0] 	       mul_out_366;
   wire [7:0] 	       mul_out_367;
   wire [7:0] 	       mul_out_368;
   wire [7:0] 	       mul_out_369;
   wire [7:0] 	       mul_out_370;
   wire [7:0] 	       mul_out_371;
   wire [7:0] 	       mul_out_372;
   wire [7:0] 	       mul_out_373;
   wire [7:0] 	       mul_out_374;
   wire [7:0] 	       mul_out_375;
   wire [7:0] 	       mul_out_376;
   wire [7:0] 	       mul_out_377;
   wire [7:0] 	       mul_out_378;
   wire [7:0] 	       mul_out_379;
   wire [7:0] 	       mul_out_380;
   wire [7:0] 	       mul_out_381;
   wire [7:0] 	       mul_out_382;
   wire [7:0] 	       mul_out_383;
   wire [7:0] 	       mul_out_384;
   wire [7:0] 	       mul_out_385;
   wire [7:0] 	       mul_out_386;
   wire [7:0] 	       mul_out_387;
   wire [7:0] 	       mul_out_388;
   wire [7:0] 	       mul_out_389;
   wire [7:0] 	       mul_out_390;
   wire [7:0] 	       mul_out_391;
   wire [7:0] 	       mul_out_392;
   wire [7:0] 	       mul_out_393;
   wire [7:0] 	       mul_out_394;
   wire [7:0] 	       mul_out_395;
   wire [7:0] 	       mul_out_396;
   wire [7:0] 	       mul_out_397;
   wire [7:0] 	       mul_out_398;
   wire [7:0] 	       mul_out_399;
   wire [7:0] 	       mul_out_400;
   wire [7:0] 	       mul_out_401;
   wire [7:0] 	       mul_out_402;
   wire [7:0] 	       mul_out_403;
   wire [7:0] 	       mul_out_404;
   wire [7:0] 	       mul_out_405;
   wire [7:0] 	       mul_out_406;
   wire [7:0] 	       mul_out_407;
   wire [7:0] 	       mul_out_408;
   wire [7:0] 	       mul_out_409;
   wire [7:0] 	       mul_out_410;
   wire [7:0] 	       mul_out_411;
   wire [7:0] 	       mul_out_412;
   wire [7:0] 	       mul_out_413;
   wire [7:0] 	       mul_out_414;
   wire [7:0] 	       mul_out_415;
   wire [7:0] 	       mul_out_416;
   wire [7:0] 	       mul_out_417;
   wire [7:0] 	       mul_out_418;
   wire [7:0] 	       mul_out_419;
   wire [7:0] 	       mul_out_420;
   wire [7:0] 	       mul_out_421;
   wire [7:0] 	       mul_out_422;
   wire [7:0] 	       mul_out_423;
   wire [7:0] 	       mul_out_424;
   wire [7:0] 	       mul_out_425;
   wire [7:0] 	       mul_out_426;
   wire [7:0] 	       mul_out_427;
   wire [7:0] 	       mul_out_428;
   wire [7:0] 	       mul_out_429;
   wire [7:0] 	       mul_out_430;
   wire [7:0] 	       mul_out_431;
   wire [7:0] 	       mul_out_432;
   wire [7:0] 	       mul_out_433;
   wire [7:0] 	       mul_out_434;
   wire [7:0] 	       mul_out_435;
   wire [7:0] 	       mul_out_436;
   wire [7:0] 	       mul_out_437;
   wire [7:0] 	       mul_out_438;
   wire [7:0] 	       mul_out_439;
   wire [7:0] 	       mul_out_440;
   wire [7:0] 	       mul_out_441;
   wire [7:0] 	       mul_out_442;
   wire [7:0] 	       mul_out_443;
   wire [7:0] 	       mul_out_444;
   wire [7:0] 	       mul_out_445;
   wire [7:0] 	       mul_out_446;
   wire [7:0] 	       mul_out_447;
   wire [7:0] 	       mul_out_448;
   wire [7:0] 	       mul_out_449;
   wire [7:0] 	       mul_out_450;
   wire [7:0] 	       mul_out_451;
   wire [7:0] 	       mul_out_452;
   wire [7:0] 	       mul_out_453;
   wire [7:0] 	       mul_out_454;
   wire [7:0] 	       mul_out_455;
   wire [7:0] 	       mul_out_456;
   wire [7:0] 	       mul_out_457;
   wire [7:0] 	       mul_out_458;
   wire [7:0] 	       mul_out_459;
   wire [7:0] 	       mul_out_460;
   wire [7:0] 	       mul_out_461;
   wire [7:0] 	       mul_out_462;
   wire [7:0] 	       mul_out_463;
   wire [7:0] 	       mul_out_464;
   wire [7:0] 	       mul_out_465;
   wire [7:0] 	       mul_out_466;
   wire [7:0] 	       mul_out_467;
   wire [7:0] 	       mul_out_468;
   wire [7:0] 	       mul_out_469;
   wire [7:0] 	       mul_out_470;
   wire [7:0] 	       mul_out_471;
   wire [7:0] 	       mul_out_472;
   wire [7:0] 	       mul_out_473;
   wire [7:0] 	       mul_out_474;
   wire [7:0] 	       mul_out_475;
   wire [7:0] 	       mul_out_476;
   wire [7:0] 	       mul_out_477;
   wire [7:0] 	       mul_out_478;
   wire [7:0] 	       mul_out_479;
   wire [7:0] 	       mul_out_480;
   wire [7:0] 	       mul_out_481;
   wire [7:0] 	       mul_out_482;
   wire [7:0] 	       mul_out_483;
   wire [7:0] 	       mul_out_484;
   wire [7:0] 	       mul_out_485;
   wire [7:0] 	       mul_out_486;
   wire [7:0] 	       mul_out_487;
   wire [7:0] 	       mul_out_488;
   wire [7:0] 	       mul_out_489;
   wire [7:0] 	       mul_out_490;
   wire [7:0] 	       mul_out_491;
   wire [7:0] 	       mul_out_492;
   wire [7:0] 	       mul_out_493;
   wire [7:0] 	       mul_out_494;
   wire [7:0] 	       mul_out_495;
   wire [7:0] 	       mul_out_496;
   wire [7:0] 	       mul_out_497;
   wire [7:0] 	       mul_out_498;
   wire [7:0] 	       mul_out_499;
   wire [7:0] 	       mul_out_500;
   wire [7:0] 	       mul_out_501;
   wire [7:0] 	       mul_out_502;
   wire [7:0] 	       mul_out_503;
   wire [7:0] 	       mul_out_504;
   wire [7:0] 	       mul_out_505;
   wire [7:0] 	       mul_out_506;
   wire [7:0] 	       mul_out_507;
   wire [7:0] 	       mul_out_508;
   wire [7:0] 	       mul_out_509;
   wire [7:0] 	       mul_out_510;
   wire [7:0] 	       mul_out_511;
   wire [7:0] 	       mul_out_512;
   wire [7:0] 	       mul_out_513;
   wire [7:0] 	       mul_out_514;
   wire [7:0] 	       mul_out_515;
   wire [7:0] 	       mul_out_516;
   wire [7:0] 	       mul_out_517;
   wire [7:0] 	       mul_out_518;
   wire [7:0] 	       mul_out_519;
   wire [7:0] 	       mul_out_520;
   wire [7:0] 	       mul_out_521;
   wire [7:0] 	       mul_out_522;
   wire [7:0] 	       mul_out_523;
   wire [7:0] 	       mul_out_524;
   wire [7:0] 	       mul_out_525;
   wire [7:0] 	       mul_out_526;
   wire [7:0] 	       mul_out_527;
   wire [7:0] 	       mul_out_528;
   wire [7:0] 	       mul_out_529;
   wire [7:0] 	       mul_out_530;
   wire [7:0] 	       mul_out_531;
   wire [7:0] 	       mul_out_532;
   wire [7:0] 	       mul_out_533;
   wire [7:0] 	       mul_out_534;
   wire [7:0] 	       mul_out_535;
   wire [7:0] 	       mul_out_536;
   wire [7:0] 	       mul_out_537;
   wire [7:0] 	       mul_out_538;
   wire [7:0] 	       mul_out_539;
   wire [7:0] 	       mul_out_540;
   wire [7:0] 	       mul_out_541;
   wire [7:0] 	       mul_out_542;
   wire [7:0] 	       mul_out_543;
   wire [7:0] 	       mul_out_544;
   wire [7:0] 	       mul_out_545;
   wire [7:0] 	       mul_out_546;
   wire [7:0] 	       mul_out_547;
   wire [7:0] 	       mul_out_548;
   wire [7:0] 	       mul_out_549;
   wire [7:0] 	       mul_out_550;
   wire [7:0] 	       mul_out_551;
   wire [7:0] 	       mul_out_552;
   wire [7:0] 	       mul_out_553;
   wire [7:0] 	       mul_out_554;
   wire [7:0] 	       mul_out_555;
   wire [7:0] 	       mul_out_556;
   wire [7:0] 	       mul_out_557;
   wire [7:0] 	       mul_out_558;
   wire [7:0] 	       mul_out_559;
   wire [7:0] 	       mul_out_560;
   wire [7:0] 	       mul_out_561;
   wire [7:0] 	       mul_out_562;
   wire [7:0] 	       mul_out_563;
   wire [7:0] 	       mul_out_564;
   wire [7:0] 	       mul_out_565;
   wire [7:0] 	       mul_out_566;
   wire [7:0] 	       mul_out_567;
   wire [7:0] 	       mul_out_568;
   wire [7:0] 	       mul_out_569;
   wire [7:0] 	       mul_out_570;
   wire [7:0] 	       mul_out_571;
   wire [7:0] 	       mul_out_572;
   wire [7:0] 	       mul_out_573;
   wire [7:0] 	       mul_out_574;
   wire [7:0] 	       mul_out_575;
   wire [7:0] 	       mul_out_576;
   wire [7:0] 	       mul_out_577;
   wire [7:0] 	       mul_out_578;
   wire [7:0] 	       mul_out_579;
   wire [7:0] 	       mul_out_580;
   wire [7:0] 	       mul_out_581;
   wire [7:0] 	       mul_out_582;
   wire [7:0] 	       mul_out_583;
   wire [7:0] 	       mul_out_584;
   wire [7:0] 	       mul_out_585;
   wire [7:0] 	       mul_out_586;
   wire [7:0] 	       mul_out_587;
   wire [7:0] 	       mul_out_588;
   wire [7:0] 	       mul_out_589;
   wire [7:0] 	       mul_out_590;
   wire [7:0] 	       mul_out_591;
   wire [7:0] 	       mul_out_592;
   wire [7:0] 	       mul_out_593;
   wire [7:0] 	       mul_out_594;
   wire [7:0] 	       mul_out_595;
   wire [7:0] 	       mul_out_596;
   wire [7:0] 	       mul_out_597;
   wire [7:0] 	       mul_out_598;
   wire [7:0] 	       mul_out_599;
   wire [7:0] 	       mul_out_600;
   wire [7:0] 	       mul_out_601;
   wire [7:0] 	       mul_out_602;
   wire [7:0] 	       mul_out_603;
   wire [7:0] 	       mul_out_604;
   wire [7:0] 	       mul_out_605;
   wire [7:0] 	       mul_out_606;
   wire [7:0] 	       mul_out_607;
   wire [7:0] 	       mul_out_608;
   wire [7:0] 	       mul_out_609;
   wire [7:0] 	       mul_out_610;
   wire [7:0] 	       mul_out_611;
   wire [7:0] 	       mul_out_612;
   wire [7:0] 	       mul_out_613;
   wire [7:0] 	       mul_out_614;
   wire [7:0] 	       mul_out_615;
   wire [7:0] 	       mul_out_616;
   wire [7:0] 	       mul_out_617;
   wire [7:0] 	       mul_out_618;
   wire [7:0] 	       mul_out_619;
   wire [7:0] 	       mul_out_620;
   wire [7:0] 	       mul_out_621;
   wire [7:0] 	       mul_out_622;
   wire [7:0] 	       mul_out_623;
   wire [7:0] 	       mul_out_624;
   wire [7:0] 	       mul_out_625;
   wire [7:0] 	       mul_out_626;
   wire [7:0] 	       mul_out_627;
   wire [7:0] 	       mul_out_628;
   wire [7:0] 	       mul_out_629;
   wire [7:0] 	       mul_out_630;
   wire [7:0] 	       mul_out_631;
   wire [7:0] 	       mul_out_632;
   wire [7:0] 	       mul_out_633;
   wire [7:0] 	       mul_out_634;
   wire [7:0] 	       mul_out_635;
   wire [7:0] 	       mul_out_636;
   wire [7:0] 	       mul_out_637;
   wire [7:0] 	       mul_out_638;
   wire [7:0] 	       mul_out_639;
   wire [7:0] 	       mul_out_640;
   wire [7:0] 	       mul_out_641;
   wire [7:0] 	       mul_out_642;
   wire [7:0] 	       mul_out_643;
   wire [7:0] 	       mul_out_644;
   wire [7:0] 	       mul_out_645;
   wire [7:0] 	       mul_out_646;
   wire [7:0] 	       mul_out_647;
   wire [7:0] 	       mul_out_648;
   wire [7:0] 	       mul_out_649;
   wire [7:0] 	       mul_out_650;
   wire [7:0] 	       mul_out_651;
   wire [7:0] 	       mul_out_652;
   wire [7:0] 	       mul_out_653;
   wire [7:0] 	       mul_out_654;
   wire [7:0] 	       mul_out_655;
   wire [7:0] 	       mul_out_656;
   wire [7:0] 	       mul_out_657;
   wire [7:0] 	       mul_out_658;
   wire [7:0] 	       mul_out_659;
   wire [7:0] 	       mul_out_660;
   wire [7:0] 	       mul_out_661;
   wire [7:0] 	       mul_out_662;
   wire [7:0] 	       mul_out_663;
   wire [7:0] 	       mul_out_664;
   wire [7:0] 	       mul_out_665;
   wire [7:0] 	       mul_out_666;
   wire [7:0] 	       mul_out_667;
   wire [7:0] 	       mul_out_668;
   wire [7:0] 	       mul_out_669;
   wire [7:0] 	       mul_out_670;
   wire [7:0] 	       mul_out_671;
   wire [7:0] 	       mul_out_672;
   wire [7:0] 	       mul_out_673;
   wire [7:0] 	       mul_out_674;
   wire [7:0] 	       mul_out_675;
   wire [7:0] 	       mul_out_676;
   wire [7:0] 	       mul_out_677;
   wire [7:0] 	       mul_out_678;
   wire [7:0] 	       mul_out_679;
   wire [7:0] 	       mul_out_680;
   wire [7:0] 	       mul_out_681;
   wire [7:0] 	       mul_out_682;
   wire [7:0] 	       mul_out_683;
   wire [7:0] 	       mul_out_684;
   wire [7:0] 	       mul_out_685;
   wire [7:0] 	       mul_out_686;
   wire [7:0] 	       mul_out_687;
   wire [7:0] 	       mul_out_688;
   wire [7:0] 	       mul_out_689;
   wire [7:0] 	       mul_out_690;
   wire [7:0] 	       mul_out_691;
   wire [7:0] 	       mul_out_692;
   wire [7:0] 	       mul_out_693;
   wire [7:0] 	       mul_out_694;
   wire [7:0] 	       mul_out_695;
   wire [7:0] 	       mul_out_696;
   wire [7:0] 	       mul_out_697;
   wire [7:0] 	       mul_out_698;
   wire [7:0] 	       mul_out_699;
   wire [7:0] 	       mul_out_700;
   wire [7:0] 	       mul_out_701;
   wire [7:0] 	       mul_out_702;
   wire [7:0] 	       mul_out_703;
   wire [7:0] 	       mul_out_704;
   wire [7:0] 	       mul_out_705;
   wire [7:0] 	       mul_out_706;
   wire [7:0] 	       mul_out_707;
   wire [7:0] 	       mul_out_708;
   wire [7:0] 	       mul_out_709;
   wire [7:0] 	       mul_out_710;
   wire [7:0] 	       mul_out_711;
   wire [7:0] 	       mul_out_712;
   wire [7:0] 	       mul_out_713;
   wire [7:0] 	       mul_out_714;
   wire [7:0] 	       mul_out_715;
   wire [7:0] 	       mul_out_716;
   wire [7:0] 	       mul_out_717;
   wire [7:0] 	       mul_out_718;
   wire [7:0] 	       mul_out_719;
   wire [7:0] 	       mul_out_720;
   wire [7:0] 	       mul_out_721;
   wire [7:0] 	       mul_out_722;
   wire [7:0] 	       mul_out_723;
   wire [7:0] 	       mul_out_724;
   wire [7:0] 	       mul_out_725;
   wire [7:0] 	       mul_out_726;
   wire [7:0] 	       mul_out_727;
   wire [7:0] 	       mul_out_728;
   wire [7:0] 	       mul_out_729;
   wire [7:0] 	       mul_out_730;
   wire [7:0] 	       mul_out_731;
   wire [7:0] 	       mul_out_732;
   wire [7:0] 	       mul_out_733;
   wire [7:0] 	       mul_out_734;
   wire [7:0] 	       mul_out_735;
   wire [7:0] 	       mul_out_736;
   wire [7:0] 	       mul_out_737;
   wire [7:0] 	       mul_out_738;
   wire [7:0] 	       mul_out_739;
   wire [7:0] 	       mul_out_740;
   wire [7:0] 	       mul_out_741;
   wire [7:0] 	       mul_out_742;
   wire [7:0] 	       mul_out_743;
   wire [7:0] 	       mul_out_744;
   wire [7:0] 	       mul_out_745;
   wire [7:0] 	       mul_out_746;
   wire [7:0] 	       mul_out_747;
   wire [7:0] 	       mul_out_748;
   wire [7:0] 	       mul_out_749;
   wire [7:0] 	       mul_out_750;
   wire [7:0] 	       mul_out_751;
   wire [7:0] 	       mul_out_752;
   wire [7:0] 	       mul_out_753;
   wire [7:0] 	       mul_out_754;
   wire [7:0] 	       mul_out_755;
   wire [7:0] 	       mul_out_756;
   wire [7:0] 	       mul_out_757;
   wire [7:0] 	       mul_out_758;
   wire [7:0] 	       mul_out_759;
   wire [7:0] 	       mul_out_760;
   wire [7:0] 	       mul_out_761;
   wire [7:0] 	       mul_out_762;
   wire [7:0] 	       mul_out_763;
   wire [7:0] 	       mul_out_764;
   wire [7:0] 	       mul_out_765;
   wire [7:0] 	       mul_out_766;
   wire [7:0] 	       mul_out_767;
   wire [7:0] 	       mul_out_768;
   wire [7:0] 	       mul_out_769;
   wire [7:0] 	       mul_out_770;
   wire [7:0] 	       mul_out_771;
   wire [7:0] 	       mul_out_772;
   wire [7:0] 	       mul_out_773;
   wire [7:0] 	       mul_out_774;
   wire [7:0] 	       mul_out_775;
   wire [7:0] 	       mul_out_776;
   wire [7:0] 	       mul_out_777;
   wire [7:0] 	       mul_out_778;
   wire [7:0] 	       mul_out_779;
   wire [7:0] 	       mul_out_780;
   wire [7:0] 	       mul_out_781;
   wire [7:0] 	       mul_out_782;
   wire [7:0] 	       mul_out_783;

   reg [20:0] 	       add_00;
   reg [20:0] 	       add_01;
   reg [20:0] 	       add_02;
   reg [20:0] 	       add_03;
   reg [20:0] 	       add_04;
   reg [20:0] 	       add_05;
   reg [20:0] 	       add_06;
   reg [20:0] 	       add_07;
   reg [20:0] 	       add_08;
   reg [20:0] 	       add_09;
   reg [20:0] 	       add_10;
   reg [20:0] 	       add_11;
   reg [20:0] 	       add_12;
   reg [20:0] 	       add_13;
   reg [20:0] 	       add_14;
   reg [20:0] 	       add_15;
   reg [20:0] 	       add_16;
   reg [20:0] 	       add_17;
   reg [20:0] 	       add_18;
   reg [20:0] 	       add_19;
   reg [20:0] 	       add_20;
   reg [20:0] 	       add_21;
   reg [20:0] 	       add_22;
   reg [20:0] 	       add_23;
   reg [20:0] 	       add_24;
   reg [20:0] 	       add_25;
   reg [20:0] 	       add_26;
   reg [20:0] 	       add_27;

   mul8x8_wrap mul_0(.CLK(CLK), .W(W[7:0]), .IMG(IMG[7:0]), .P(mul_out_0));
   mul8x8_wrap mul_1(.CLK(CLK), .W(W[15:8]), .IMG(IMG[15:8]), .P(mul_out_1));
   mul8x8_wrap mul_2(.CLK(CLK), .W(W[23:16]), .IMG(IMG[23:16]), .P(mul_out_2));
   mul8x8_wrap mul_3(.CLK(CLK), .W(W[31:24]), .IMG(IMG[31:24]), .P(mul_out_3));
   mul8x8_wrap mul_4(.CLK(CLK), .W(W[39:32]), .IMG(IMG[39:32]), .P(mul_out_4));
   mul8x8_wrap mul_5(.CLK(CLK), .W(W[47:40]), .IMG(IMG[47:40]), .P(mul_out_5));
   mul8x8_wrap mul_6(.CLK(CLK), .W(W[55:48]), .IMG(IMG[55:48]), .P(mul_out_6));
   mul8x8_wrap mul_7(.CLK(CLK), .W(W[63:56]), .IMG(IMG[63:56]), .P(mul_out_7));
   mul8x8_wrap mul_8(.CLK(CLK), .W(W[71:64]), .IMG(IMG[71:64]), .P(mul_out_8));
   mul8x8_wrap mul_9(.CLK(CLK), .W(W[79:72]), .IMG(IMG[79:72]), .P(mul_out_9));
   mul8x8_wrap mul_10(.CLK(CLK), .W(W[87:80]), .IMG(IMG[87:80]), .P(mul_out_10));
   mul8x8_wrap mul_11(.CLK(CLK), .W(W[95:88]), .IMG(IMG[95:88]), .P(mul_out_11));
   mul8x8_wrap mul_12(.CLK(CLK), .W(W[103:96]), .IMG(IMG[103:96]), .P(mul_out_12));
   mul8x8_wrap mul_13(.CLK(CLK), .W(W[111:104]), .IMG(IMG[111:104]), .P(mul_out_13));
   mul8x8_wrap mul_14(.CLK(CLK), .W(W[119:112]), .IMG(IMG[119:112]), .P(mul_out_14));
   mul8x8_wrap mul_15(.CLK(CLK), .W(W[127:120]), .IMG(IMG[127:120]), .P(mul_out_15));
   mul8x8_wrap mul_16(.CLK(CLK), .W(W[135:128]), .IMG(IMG[135:128]), .P(mul_out_16));
   mul8x8_wrap mul_17(.CLK(CLK), .W(W[143:136]), .IMG(IMG[143:136]), .P(mul_out_17));
   mul8x8_wrap mul_18(.CLK(CLK), .W(W[151:144]), .IMG(IMG[151:144]), .P(mul_out_18));
   mul8x8_wrap mul_19(.CLK(CLK), .W(W[159:152]), .IMG(IMG[159:152]), .P(mul_out_19));
   mul8x8_wrap mul_20(.CLK(CLK), .W(W[167:160]), .IMG(IMG[167:160]), .P(mul_out_20));
   mul8x8_wrap mul_21(.CLK(CLK), .W(W[175:168]), .IMG(IMG[175:168]), .P(mul_out_21));
   mul8x8_wrap mul_22(.CLK(CLK), .W(W[183:176]), .IMG(IMG[183:176]), .P(mul_out_22));
   mul8x8_wrap mul_23(.CLK(CLK), .W(W[191:184]), .IMG(IMG[191:184]), .P(mul_out_23));
   mul8x8_wrap mul_24(.CLK(CLK), .W(W[199:192]), .IMG(IMG[199:192]), .P(mul_out_24));
   mul8x8_wrap mul_25(.CLK(CLK), .W(W[207:200]), .IMG(IMG[207:200]), .P(mul_out_25));
   mul8x8_wrap mul_26(.CLK(CLK), .W(W[215:208]), .IMG(IMG[215:208]), .P(mul_out_26));
   mul8x8_wrap mul_27(.CLK(CLK), .W(W[223:216]), .IMG(IMG[223:216]), .P(mul_out_27));
   mul8x8_wrap mul_28(.CLK(CLK), .W(W[231:224]), .IMG(IMG[231:224]), .P(mul_out_28));
   mul8x8_wrap mul_29(.CLK(CLK), .W(W[239:232]), .IMG(IMG[239:232]), .P(mul_out_29));
   mul8x8_wrap mul_30(.CLK(CLK), .W(W[247:240]), .IMG(IMG[247:240]), .P(mul_out_30));
   mul8x8_wrap mul_31(.CLK(CLK), .W(W[255:248]), .IMG(IMG[255:248]), .P(mul_out_31));
   mul8x8_wrap mul_32(.CLK(CLK), .W(W[263:256]), .IMG(IMG[263:256]), .P(mul_out_32));
   mul8x8_wrap mul_33(.CLK(CLK), .W(W[271:264]), .IMG(IMG[271:264]), .P(mul_out_33));
   mul8x8_wrap mul_34(.CLK(CLK), .W(W[279:272]), .IMG(IMG[279:272]), .P(mul_out_34));
   mul8x8_wrap mul_35(.CLK(CLK), .W(W[287:280]), .IMG(IMG[287:280]), .P(mul_out_35));
   mul8x8_wrap mul_36(.CLK(CLK), .W(W[295:288]), .IMG(IMG[295:288]), .P(mul_out_36));
   mul8x8_wrap mul_37(.CLK(CLK), .W(W[303:296]), .IMG(IMG[303:296]), .P(mul_out_37));
   mul8x8_wrap mul_38(.CLK(CLK), .W(W[311:304]), .IMG(IMG[311:304]), .P(mul_out_38));
   mul8x8_wrap mul_39(.CLK(CLK), .W(W[319:312]), .IMG(IMG[319:312]), .P(mul_out_39));
   mul8x8_wrap mul_40(.CLK(CLK), .W(W[327:320]), .IMG(IMG[327:320]), .P(mul_out_40));
   mul8x8_wrap mul_41(.CLK(CLK), .W(W[335:328]), .IMG(IMG[335:328]), .P(mul_out_41));
   mul8x8_wrap mul_42(.CLK(CLK), .W(W[343:336]), .IMG(IMG[343:336]), .P(mul_out_42));
   mul8x8_wrap mul_43(.CLK(CLK), .W(W[351:344]), .IMG(IMG[351:344]), .P(mul_out_43));
   mul8x8_wrap mul_44(.CLK(CLK), .W(W[359:352]), .IMG(IMG[359:352]), .P(mul_out_44));
   mul8x8_wrap mul_45(.CLK(CLK), .W(W[367:360]), .IMG(IMG[367:360]), .P(mul_out_45));
   mul8x8_wrap mul_46(.CLK(CLK), .W(W[375:368]), .IMG(IMG[375:368]), .P(mul_out_46));
   mul8x8_wrap mul_47(.CLK(CLK), .W(W[383:376]), .IMG(IMG[383:376]), .P(mul_out_47));
   mul8x8_wrap mul_48(.CLK(CLK), .W(W[391:384]), .IMG(IMG[391:384]), .P(mul_out_48));
   mul8x8_wrap mul_49(.CLK(CLK), .W(W[399:392]), .IMG(IMG[399:392]), .P(mul_out_49));
   mul8x8_wrap mul_50(.CLK(CLK), .W(W[407:400]), .IMG(IMG[407:400]), .P(mul_out_50));
   mul8x8_wrap mul_51(.CLK(CLK), .W(W[415:408]), .IMG(IMG[415:408]), .P(mul_out_51));
   mul8x8_wrap mul_52(.CLK(CLK), .W(W[423:416]), .IMG(IMG[423:416]), .P(mul_out_52));
   mul8x8_wrap mul_53(.CLK(CLK), .W(W[431:424]), .IMG(IMG[431:424]), .P(mul_out_53));
   mul8x8_wrap mul_54(.CLK(CLK), .W(W[439:432]), .IMG(IMG[439:432]), .P(mul_out_54));
   mul8x8_wrap mul_55(.CLK(CLK), .W(W[447:440]), .IMG(IMG[447:440]), .P(mul_out_55));
   mul8x8_wrap mul_56(.CLK(CLK), .W(W[455:448]), .IMG(IMG[455:448]), .P(mul_out_56));
   mul8x8_wrap mul_57(.CLK(CLK), .W(W[463:456]), .IMG(IMG[463:456]), .P(mul_out_57));
   mul8x8_wrap mul_58(.CLK(CLK), .W(W[471:464]), .IMG(IMG[471:464]), .P(mul_out_58));
   mul8x8_wrap mul_59(.CLK(CLK), .W(W[479:472]), .IMG(IMG[479:472]), .P(mul_out_59));
   mul8x8_wrap mul_60(.CLK(CLK), .W(W[487:480]), .IMG(IMG[487:480]), .P(mul_out_60));
   mul8x8_wrap mul_61(.CLK(CLK), .W(W[495:488]), .IMG(IMG[495:488]), .P(mul_out_61));
   mul8x8_wrap mul_62(.CLK(CLK), .W(W[503:496]), .IMG(IMG[503:496]), .P(mul_out_62));
   mul8x8_wrap mul_63(.CLK(CLK), .W(W[511:504]), .IMG(IMG[511:504]), .P(mul_out_63));
   mul8x8_wrap mul_64(.CLK(CLK), .W(W[519:512]), .IMG(IMG[519:512]), .P(mul_out_64));
   mul8x8_wrap mul_65(.CLK(CLK), .W(W[527:520]), .IMG(IMG[527:520]), .P(mul_out_65));
   mul8x8_wrap mul_66(.CLK(CLK), .W(W[535:528]), .IMG(IMG[535:528]), .P(mul_out_66));
   mul8x8_wrap mul_67(.CLK(CLK), .W(W[543:536]), .IMG(IMG[543:536]), .P(mul_out_67));
   mul8x8_wrap mul_68(.CLK(CLK), .W(W[551:544]), .IMG(IMG[551:544]), .P(mul_out_68));
   mul8x8_wrap mul_69(.CLK(CLK), .W(W[559:552]), .IMG(IMG[559:552]), .P(mul_out_69));
   mul8x8_wrap mul_70(.CLK(CLK), .W(W[567:560]), .IMG(IMG[567:560]), .P(mul_out_70));
   mul8x8_wrap mul_71(.CLK(CLK), .W(W[575:568]), .IMG(IMG[575:568]), .P(mul_out_71));
   mul8x8_wrap mul_72(.CLK(CLK), .W(W[583:576]), .IMG(IMG[583:576]), .P(mul_out_72));
   mul8x8_wrap mul_73(.CLK(CLK), .W(W[591:584]), .IMG(IMG[591:584]), .P(mul_out_73));
   mul8x8_wrap mul_74(.CLK(CLK), .W(W[599:592]), .IMG(IMG[599:592]), .P(mul_out_74));
   mul8x8_wrap mul_75(.CLK(CLK), .W(W[607:600]), .IMG(IMG[607:600]), .P(mul_out_75));
   mul8x8_wrap mul_76(.CLK(CLK), .W(W[615:608]), .IMG(IMG[615:608]), .P(mul_out_76));
   mul8x8_wrap mul_77(.CLK(CLK), .W(W[623:616]), .IMG(IMG[623:616]), .P(mul_out_77));
   mul8x8_wrap mul_78(.CLK(CLK), .W(W[631:624]), .IMG(IMG[631:624]), .P(mul_out_78));
   mul8x8_wrap mul_79(.CLK(CLK), .W(W[639:632]), .IMG(IMG[639:632]), .P(mul_out_79));
   mul8x8_wrap mul_80(.CLK(CLK), .W(W[647:640]), .IMG(IMG[647:640]), .P(mul_out_80));
   mul8x8_wrap mul_81(.CLK(CLK), .W(W[655:648]), .IMG(IMG[655:648]), .P(mul_out_81));
   mul8x8_wrap mul_82(.CLK(CLK), .W(W[663:656]), .IMG(IMG[663:656]), .P(mul_out_82));
   mul8x8_wrap mul_83(.CLK(CLK), .W(W[671:664]), .IMG(IMG[671:664]), .P(mul_out_83));
   mul8x8_wrap mul_84(.CLK(CLK), .W(W[679:672]), .IMG(IMG[679:672]), .P(mul_out_84));
   mul8x8_wrap mul_85(.CLK(CLK), .W(W[687:680]), .IMG(IMG[687:680]), .P(mul_out_85));
   mul8x8_wrap mul_86(.CLK(CLK), .W(W[695:688]), .IMG(IMG[695:688]), .P(mul_out_86));
   mul8x8_wrap mul_87(.CLK(CLK), .W(W[703:696]), .IMG(IMG[703:696]), .P(mul_out_87));
   mul8x8_wrap mul_88(.CLK(CLK), .W(W[711:704]), .IMG(IMG[711:704]), .P(mul_out_88));
   mul8x8_wrap mul_89(.CLK(CLK), .W(W[719:712]), .IMG(IMG[719:712]), .P(mul_out_89));
   mul8x8_wrap mul_90(.CLK(CLK), .W(W[727:720]), .IMG(IMG[727:720]), .P(mul_out_90));
   mul8x8_wrap mul_91(.CLK(CLK), .W(W[735:728]), .IMG(IMG[735:728]), .P(mul_out_91));
   mul8x8_wrap mul_92(.CLK(CLK), .W(W[743:736]), .IMG(IMG[743:736]), .P(mul_out_92));
   mul8x8_wrap mul_93(.CLK(CLK), .W(W[751:744]), .IMG(IMG[751:744]), .P(mul_out_93));
   mul8x8_wrap mul_94(.CLK(CLK), .W(W[759:752]), .IMG(IMG[759:752]), .P(mul_out_94));
   mul8x8_wrap mul_95(.CLK(CLK), .W(W[767:760]), .IMG(IMG[767:760]), .P(mul_out_95));
   mul8x8_wrap mul_96(.CLK(CLK), .W(W[775:768]), .IMG(IMG[775:768]), .P(mul_out_96));
   mul8x8_wrap mul_97(.CLK(CLK), .W(W[783:776]), .IMG(IMG[783:776]), .P(mul_out_97));
   mul8x8_wrap mul_98(.CLK(CLK), .W(W[791:784]), .IMG(IMG[791:784]), .P(mul_out_98));
   mul8x8_wrap mul_99(.CLK(CLK), .W(W[799:792]), .IMG(IMG[799:792]), .P(mul_out_99));
   mul8x8_wrap mul_100(.CLK(CLK), .W(W[807:800]), .IMG(IMG[807:800]), .P(mul_out_100));
   mul8x8_wrap mul_101(.CLK(CLK), .W(W[815:808]), .IMG(IMG[815:808]), .P(mul_out_101));
   mul8x8_wrap mul_102(.CLK(CLK), .W(W[823:816]), .IMG(IMG[823:816]), .P(mul_out_102));
   mul8x8_wrap mul_103(.CLK(CLK), .W(W[831:824]), .IMG(IMG[831:824]), .P(mul_out_103));
   mul8x8_wrap mul_104(.CLK(CLK), .W(W[839:832]), .IMG(IMG[839:832]), .P(mul_out_104));
   mul8x8_wrap mul_105(.CLK(CLK), .W(W[847:840]), .IMG(IMG[847:840]), .P(mul_out_105));
   mul8x8_wrap mul_106(.CLK(CLK), .W(W[855:848]), .IMG(IMG[855:848]), .P(mul_out_106));
   mul8x8_wrap mul_107(.CLK(CLK), .W(W[863:856]), .IMG(IMG[863:856]), .P(mul_out_107));
   mul8x8_wrap mul_108(.CLK(CLK), .W(W[871:864]), .IMG(IMG[871:864]), .P(mul_out_108));
   mul8x8_wrap mul_109(.CLK(CLK), .W(W[879:872]), .IMG(IMG[879:872]), .P(mul_out_109));
   mul8x8_wrap mul_110(.CLK(CLK), .W(W[887:880]), .IMG(IMG[887:880]), .P(mul_out_110));
   mul8x8_wrap mul_111(.CLK(CLK), .W(W[895:888]), .IMG(IMG[895:888]), .P(mul_out_111));
   mul8x8_wrap mul_112(.CLK(CLK), .W(W[903:896]), .IMG(IMG[903:896]), .P(mul_out_112));
   mul8x8_wrap mul_113(.CLK(CLK), .W(W[911:904]), .IMG(IMG[911:904]), .P(mul_out_113));
   mul8x8_wrap mul_114(.CLK(CLK), .W(W[919:912]), .IMG(IMG[919:912]), .P(mul_out_114));
   mul8x8_wrap mul_115(.CLK(CLK), .W(W[927:920]), .IMG(IMG[927:920]), .P(mul_out_115));
   mul8x8_wrap mul_116(.CLK(CLK), .W(W[935:928]), .IMG(IMG[935:928]), .P(mul_out_116));
   mul8x8_wrap mul_117(.CLK(CLK), .W(W[943:936]), .IMG(IMG[943:936]), .P(mul_out_117));
   mul8x8_wrap mul_118(.CLK(CLK), .W(W[951:944]), .IMG(IMG[951:944]), .P(mul_out_118));
   mul8x8_wrap mul_119(.CLK(CLK), .W(W[959:952]), .IMG(IMG[959:952]), .P(mul_out_119));
   mul8x8_wrap mul_120(.CLK(CLK), .W(W[967:960]), .IMG(IMG[967:960]), .P(mul_out_120));
   mul8x8_wrap mul_121(.CLK(CLK), .W(W[975:968]), .IMG(IMG[975:968]), .P(mul_out_121));
   mul8x8_wrap mul_122(.CLK(CLK), .W(W[983:976]), .IMG(IMG[983:976]), .P(mul_out_122));
   mul8x8_wrap mul_123(.CLK(CLK), .W(W[991:984]), .IMG(IMG[991:984]), .P(mul_out_123));
   mul8x8_wrap mul_124(.CLK(CLK), .W(W[999:992]), .IMG(IMG[999:992]), .P(mul_out_124));
   mul8x8_wrap mul_125(.CLK(CLK), .W(W[1007:1000]), .IMG(IMG[1007:1000]), .P(mul_out_125));
   mul8x8_wrap mul_126(.CLK(CLK), .W(W[1015:1008]), .IMG(IMG[1015:1008]), .P(mul_out_126));
   mul8x8_wrap mul_127(.CLK(CLK), .W(W[1023:1016]), .IMG(IMG[1023:1016]), .P(mul_out_127));
   mul8x8_wrap mul_128(.CLK(CLK), .W(W[1031:1024]), .IMG(IMG[1031:1024]), .P(mul_out_128));
   mul8x8_wrap mul_129(.CLK(CLK), .W(W[1039:1032]), .IMG(IMG[1039:1032]), .P(mul_out_129));
   mul8x8_wrap mul_130(.CLK(CLK), .W(W[1047:1040]), .IMG(IMG[1047:1040]), .P(mul_out_130));
   mul8x8_wrap mul_131(.CLK(CLK), .W(W[1055:1048]), .IMG(IMG[1055:1048]), .P(mul_out_131));
   mul8x8_wrap mul_132(.CLK(CLK), .W(W[1063:1056]), .IMG(IMG[1063:1056]), .P(mul_out_132));
   mul8x8_wrap mul_133(.CLK(CLK), .W(W[1071:1064]), .IMG(IMG[1071:1064]), .P(mul_out_133));
   mul8x8_wrap mul_134(.CLK(CLK), .W(W[1079:1072]), .IMG(IMG[1079:1072]), .P(mul_out_134));
   mul8x8_wrap mul_135(.CLK(CLK), .W(W[1087:1080]), .IMG(IMG[1087:1080]), .P(mul_out_135));
   mul8x8_wrap mul_136(.CLK(CLK), .W(W[1095:1088]), .IMG(IMG[1095:1088]), .P(mul_out_136));
   mul8x8_wrap mul_137(.CLK(CLK), .W(W[1103:1096]), .IMG(IMG[1103:1096]), .P(mul_out_137));
   mul8x8_wrap mul_138(.CLK(CLK), .W(W[1111:1104]), .IMG(IMG[1111:1104]), .P(mul_out_138));
   mul8x8_wrap mul_139(.CLK(CLK), .W(W[1119:1112]), .IMG(IMG[1119:1112]), .P(mul_out_139));
   mul8x8_wrap mul_140(.CLK(CLK), .W(W[1127:1120]), .IMG(IMG[1127:1120]), .P(mul_out_140));
   mul8x8_wrap mul_141(.CLK(CLK), .W(W[1135:1128]), .IMG(IMG[1135:1128]), .P(mul_out_141));
   mul8x8_wrap mul_142(.CLK(CLK), .W(W[1143:1136]), .IMG(IMG[1143:1136]), .P(mul_out_142));
   mul8x8_wrap mul_143(.CLK(CLK), .W(W[1151:1144]), .IMG(IMG[1151:1144]), .P(mul_out_143));
   mul8x8_wrap mul_144(.CLK(CLK), .W(W[1159:1152]), .IMG(IMG[1159:1152]), .P(mul_out_144));
   mul8x8_wrap mul_145(.CLK(CLK), .W(W[1167:1160]), .IMG(IMG[1167:1160]), .P(mul_out_145));
   mul8x8_wrap mul_146(.CLK(CLK), .W(W[1175:1168]), .IMG(IMG[1175:1168]), .P(mul_out_146));
   mul8x8_wrap mul_147(.CLK(CLK), .W(W[1183:1176]), .IMG(IMG[1183:1176]), .P(mul_out_147));
   mul8x8_wrap mul_148(.CLK(CLK), .W(W[1191:1184]), .IMG(IMG[1191:1184]), .P(mul_out_148));
   mul8x8_wrap mul_149(.CLK(CLK), .W(W[1199:1192]), .IMG(IMG[1199:1192]), .P(mul_out_149));
   mul8x8_wrap mul_150(.CLK(CLK), .W(W[1207:1200]), .IMG(IMG[1207:1200]), .P(mul_out_150));
   mul8x8_wrap mul_151(.CLK(CLK), .W(W[1215:1208]), .IMG(IMG[1215:1208]), .P(mul_out_151));
   mul8x8_wrap mul_152(.CLK(CLK), .W(W[1223:1216]), .IMG(IMG[1223:1216]), .P(mul_out_152));
   mul8x8_wrap mul_153(.CLK(CLK), .W(W[1231:1224]), .IMG(IMG[1231:1224]), .P(mul_out_153));
   mul8x8_wrap mul_154(.CLK(CLK), .W(W[1239:1232]), .IMG(IMG[1239:1232]), .P(mul_out_154));
   mul8x8_wrap mul_155(.CLK(CLK), .W(W[1247:1240]), .IMG(IMG[1247:1240]), .P(mul_out_155));
   mul8x8_wrap mul_156(.CLK(CLK), .W(W[1255:1248]), .IMG(IMG[1255:1248]), .P(mul_out_156));
   mul8x8_wrap mul_157(.CLK(CLK), .W(W[1263:1256]), .IMG(IMG[1263:1256]), .P(mul_out_157));
   mul8x8_wrap mul_158(.CLK(CLK), .W(W[1271:1264]), .IMG(IMG[1271:1264]), .P(mul_out_158));
   mul8x8_wrap mul_159(.CLK(CLK), .W(W[1279:1272]), .IMG(IMG[1279:1272]), .P(mul_out_159));
   mul8x8_wrap mul_160(.CLK(CLK), .W(W[1287:1280]), .IMG(IMG[1287:1280]), .P(mul_out_160));
   mul8x8_wrap mul_161(.CLK(CLK), .W(W[1295:1288]), .IMG(IMG[1295:1288]), .P(mul_out_161));
   mul8x8_wrap mul_162(.CLK(CLK), .W(W[1303:1296]), .IMG(IMG[1303:1296]), .P(mul_out_162));
   mul8x8_wrap mul_163(.CLK(CLK), .W(W[1311:1304]), .IMG(IMG[1311:1304]), .P(mul_out_163));
   mul8x8_wrap mul_164(.CLK(CLK), .W(W[1319:1312]), .IMG(IMG[1319:1312]), .P(mul_out_164));
   mul8x8_wrap mul_165(.CLK(CLK), .W(W[1327:1320]), .IMG(IMG[1327:1320]), .P(mul_out_165));
   mul8x8_wrap mul_166(.CLK(CLK), .W(W[1335:1328]), .IMG(IMG[1335:1328]), .P(mul_out_166));
   mul8x8_wrap mul_167(.CLK(CLK), .W(W[1343:1336]), .IMG(IMG[1343:1336]), .P(mul_out_167));
   mul8x8_wrap mul_168(.CLK(CLK), .W(W[1351:1344]), .IMG(IMG[1351:1344]), .P(mul_out_168));
   mul8x8_wrap mul_169(.CLK(CLK), .W(W[1359:1352]), .IMG(IMG[1359:1352]), .P(mul_out_169));
   mul8x8_wrap mul_170(.CLK(CLK), .W(W[1367:1360]), .IMG(IMG[1367:1360]), .P(mul_out_170));
   mul8x8_wrap mul_171(.CLK(CLK), .W(W[1375:1368]), .IMG(IMG[1375:1368]), .P(mul_out_171));
   mul8x8_wrap mul_172(.CLK(CLK), .W(W[1383:1376]), .IMG(IMG[1383:1376]), .P(mul_out_172));
   mul8x8_wrap mul_173(.CLK(CLK), .W(W[1391:1384]), .IMG(IMG[1391:1384]), .P(mul_out_173));
   mul8x8_wrap mul_174(.CLK(CLK), .W(W[1399:1392]), .IMG(IMG[1399:1392]), .P(mul_out_174));
   mul8x8_wrap mul_175(.CLK(CLK), .W(W[1407:1400]), .IMG(IMG[1407:1400]), .P(mul_out_175));
   mul8x8_wrap mul_176(.CLK(CLK), .W(W[1415:1408]), .IMG(IMG[1415:1408]), .P(mul_out_176));
   mul8x8_wrap mul_177(.CLK(CLK), .W(W[1423:1416]), .IMG(IMG[1423:1416]), .P(mul_out_177));
   mul8x8_wrap mul_178(.CLK(CLK), .W(W[1431:1424]), .IMG(IMG[1431:1424]), .P(mul_out_178));
   mul8x8_wrap mul_179(.CLK(CLK), .W(W[1439:1432]), .IMG(IMG[1439:1432]), .P(mul_out_179));
   mul8x8_wrap mul_180(.CLK(CLK), .W(W[1447:1440]), .IMG(IMG[1447:1440]), .P(mul_out_180));
   mul8x8_wrap mul_181(.CLK(CLK), .W(W[1455:1448]), .IMG(IMG[1455:1448]), .P(mul_out_181));
   mul8x8_wrap mul_182(.CLK(CLK), .W(W[1463:1456]), .IMG(IMG[1463:1456]), .P(mul_out_182));
   mul8x8_wrap mul_183(.CLK(CLK), .W(W[1471:1464]), .IMG(IMG[1471:1464]), .P(mul_out_183));
   mul8x8_wrap mul_184(.CLK(CLK), .W(W[1479:1472]), .IMG(IMG[1479:1472]), .P(mul_out_184));
   mul8x8_wrap mul_185(.CLK(CLK), .W(W[1487:1480]), .IMG(IMG[1487:1480]), .P(mul_out_185));
   mul8x8_wrap mul_186(.CLK(CLK), .W(W[1495:1488]), .IMG(IMG[1495:1488]), .P(mul_out_186));
   mul8x8_wrap mul_187(.CLK(CLK), .W(W[1503:1496]), .IMG(IMG[1503:1496]), .P(mul_out_187));
   mul8x8_wrap mul_188(.CLK(CLK), .W(W[1511:1504]), .IMG(IMG[1511:1504]), .P(mul_out_188));
   mul8x8_wrap mul_189(.CLK(CLK), .W(W[1519:1512]), .IMG(IMG[1519:1512]), .P(mul_out_189));
   mul8x8_wrap mul_190(.CLK(CLK), .W(W[1527:1520]), .IMG(IMG[1527:1520]), .P(mul_out_190));
   mul8x8_wrap mul_191(.CLK(CLK), .W(W[1535:1528]), .IMG(IMG[1535:1528]), .P(mul_out_191));
   mul8x8_wrap mul_192(.CLK(CLK), .W(W[1543:1536]), .IMG(IMG[1543:1536]), .P(mul_out_192));
   mul8x8_wrap mul_193(.CLK(CLK), .W(W[1551:1544]), .IMG(IMG[1551:1544]), .P(mul_out_193));
   mul8x8_wrap mul_194(.CLK(CLK), .W(W[1559:1552]), .IMG(IMG[1559:1552]), .P(mul_out_194));
   mul8x8_wrap mul_195(.CLK(CLK), .W(W[1567:1560]), .IMG(IMG[1567:1560]), .P(mul_out_195));
   mul8x8_wrap mul_196(.CLK(CLK), .W(W[1575:1568]), .IMG(IMG[1575:1568]), .P(mul_out_196));
   mul8x8_wrap mul_197(.CLK(CLK), .W(W[1583:1576]), .IMG(IMG[1583:1576]), .P(mul_out_197));
   mul8x8_wrap mul_198(.CLK(CLK), .W(W[1591:1584]), .IMG(IMG[1591:1584]), .P(mul_out_198));
   mul8x8_wrap mul_199(.CLK(CLK), .W(W[1599:1592]), .IMG(IMG[1599:1592]), .P(mul_out_199));
   mul8x8_wrap mul_200(.CLK(CLK), .W(W[1607:1600]), .IMG(IMG[1607:1600]), .P(mul_out_200));
   mul8x8_wrap mul_201(.CLK(CLK), .W(W[1615:1608]), .IMG(IMG[1615:1608]), .P(mul_out_201));
   mul8x8_wrap mul_202(.CLK(CLK), .W(W[1623:1616]), .IMG(IMG[1623:1616]), .P(mul_out_202));
   mul8x8_wrap mul_203(.CLK(CLK), .W(W[1631:1624]), .IMG(IMG[1631:1624]), .P(mul_out_203));
   mul8x8_wrap mul_204(.CLK(CLK), .W(W[1639:1632]), .IMG(IMG[1639:1632]), .P(mul_out_204));
   mul8x8_wrap mul_205(.CLK(CLK), .W(W[1647:1640]), .IMG(IMG[1647:1640]), .P(mul_out_205));
   mul8x8_wrap mul_206(.CLK(CLK), .W(W[1655:1648]), .IMG(IMG[1655:1648]), .P(mul_out_206));
   mul8x8_wrap mul_207(.CLK(CLK), .W(W[1663:1656]), .IMG(IMG[1663:1656]), .P(mul_out_207));
   mul8x8_wrap mul_208(.CLK(CLK), .W(W[1671:1664]), .IMG(IMG[1671:1664]), .P(mul_out_208));
   mul8x8_wrap mul_209(.CLK(CLK), .W(W[1679:1672]), .IMG(IMG[1679:1672]), .P(mul_out_209));
   mul8x8_wrap mul_210(.CLK(CLK), .W(W[1687:1680]), .IMG(IMG[1687:1680]), .P(mul_out_210));
   mul8x8_wrap mul_211(.CLK(CLK), .W(W[1695:1688]), .IMG(IMG[1695:1688]), .P(mul_out_211));
   mul8x8_wrap mul_212(.CLK(CLK), .W(W[1703:1696]), .IMG(IMG[1703:1696]), .P(mul_out_212));
   mul8x8_wrap mul_213(.CLK(CLK), .W(W[1711:1704]), .IMG(IMG[1711:1704]), .P(mul_out_213));
   mul8x8_wrap mul_214(.CLK(CLK), .W(W[1719:1712]), .IMG(IMG[1719:1712]), .P(mul_out_214));
   mul8x8_wrap mul_215(.CLK(CLK), .W(W[1727:1720]), .IMG(IMG[1727:1720]), .P(mul_out_215));
   mul8x8_wrap mul_216(.CLK(CLK), .W(W[1735:1728]), .IMG(IMG[1735:1728]), .P(mul_out_216));
   mul8x8_wrap mul_217(.CLK(CLK), .W(W[1743:1736]), .IMG(IMG[1743:1736]), .P(mul_out_217));
   mul8x8_wrap mul_218(.CLK(CLK), .W(W[1751:1744]), .IMG(IMG[1751:1744]), .P(mul_out_218));
   mul8x8_wrap mul_219(.CLK(CLK), .W(W[1759:1752]), .IMG(IMG[1759:1752]), .P(mul_out_219));
   mul8x8_wrap mul_220(.CLK(CLK), .W(W[1767:1760]), .IMG(IMG[1767:1760]), .P(mul_out_220));
   mul8x8_wrap mul_221(.CLK(CLK), .W(W[1775:1768]), .IMG(IMG[1775:1768]), .P(mul_out_221));
   mul8x8_wrap mul_222(.CLK(CLK), .W(W[1783:1776]), .IMG(IMG[1783:1776]), .P(mul_out_222));
   mul8x8_wrap mul_223(.CLK(CLK), .W(W[1791:1784]), .IMG(IMG[1791:1784]), .P(mul_out_223));
   mul8x8_wrap mul_224(.CLK(CLK), .W(W[1799:1792]), .IMG(IMG[1799:1792]), .P(mul_out_224));
   mul8x8_wrap mul_225(.CLK(CLK), .W(W[1807:1800]), .IMG(IMG[1807:1800]), .P(mul_out_225));
   mul8x8_wrap mul_226(.CLK(CLK), .W(W[1815:1808]), .IMG(IMG[1815:1808]), .P(mul_out_226));
   mul8x8_wrap mul_227(.CLK(CLK), .W(W[1823:1816]), .IMG(IMG[1823:1816]), .P(mul_out_227));
   mul8x8_wrap mul_228(.CLK(CLK), .W(W[1831:1824]), .IMG(IMG[1831:1824]), .P(mul_out_228));
   mul8x8_wrap mul_229(.CLK(CLK), .W(W[1839:1832]), .IMG(IMG[1839:1832]), .P(mul_out_229));
   mul8x8_wrap mul_230(.CLK(CLK), .W(W[1847:1840]), .IMG(IMG[1847:1840]), .P(mul_out_230));
   mul8x8_wrap mul_231(.CLK(CLK), .W(W[1855:1848]), .IMG(IMG[1855:1848]), .P(mul_out_231));
   mul8x8_wrap mul_232(.CLK(CLK), .W(W[1863:1856]), .IMG(IMG[1863:1856]), .P(mul_out_232));
   mul8x8_wrap mul_233(.CLK(CLK), .W(W[1871:1864]), .IMG(IMG[1871:1864]), .P(mul_out_233));
   mul8x8_wrap mul_234(.CLK(CLK), .W(W[1879:1872]), .IMG(IMG[1879:1872]), .P(mul_out_234));
   mul8x8_wrap mul_235(.CLK(CLK), .W(W[1887:1880]), .IMG(IMG[1887:1880]), .P(mul_out_235));
   mul8x8_wrap mul_236(.CLK(CLK), .W(W[1895:1888]), .IMG(IMG[1895:1888]), .P(mul_out_236));
   mul8x8_wrap mul_237(.CLK(CLK), .W(W[1903:1896]), .IMG(IMG[1903:1896]), .P(mul_out_237));
   mul8x8_wrap mul_238(.CLK(CLK), .W(W[1911:1904]), .IMG(IMG[1911:1904]), .P(mul_out_238));
   mul8x8_wrap mul_239(.CLK(CLK), .W(W[1919:1912]), .IMG(IMG[1919:1912]), .P(mul_out_239));
   mul8x8_wrap mul_240(.CLK(CLK), .W(W[1927:1920]), .IMG(IMG[1927:1920]), .P(mul_out_240));
   mul8x8_wrap mul_241(.CLK(CLK), .W(W[1935:1928]), .IMG(IMG[1935:1928]), .P(mul_out_241));
   mul8x8_wrap mul_242(.CLK(CLK), .W(W[1943:1936]), .IMG(IMG[1943:1936]), .P(mul_out_242));
   mul8x8_wrap mul_243(.CLK(CLK), .W(W[1951:1944]), .IMG(IMG[1951:1944]), .P(mul_out_243));
   mul8x8_wrap mul_244(.CLK(CLK), .W(W[1959:1952]), .IMG(IMG[1959:1952]), .P(mul_out_244));
   mul8x8_wrap mul_245(.CLK(CLK), .W(W[1967:1960]), .IMG(IMG[1967:1960]), .P(mul_out_245));
   mul8x8_wrap mul_246(.CLK(CLK), .W(W[1975:1968]), .IMG(IMG[1975:1968]), .P(mul_out_246));
   mul8x8_wrap mul_247(.CLK(CLK), .W(W[1983:1976]), .IMG(IMG[1983:1976]), .P(mul_out_247));
   mul8x8_wrap mul_248(.CLK(CLK), .W(W[1991:1984]), .IMG(IMG[1991:1984]), .P(mul_out_248));
   mul8x8_wrap mul_249(.CLK(CLK), .W(W[1999:1992]), .IMG(IMG[1999:1992]), .P(mul_out_249));
   mul8x8_wrap mul_250(.CLK(CLK), .W(W[2007:2000]), .IMG(IMG[2007:2000]), .P(mul_out_250));
   mul8x8_wrap mul_251(.CLK(CLK), .W(W[2015:2008]), .IMG(IMG[2015:2008]), .P(mul_out_251));
   mul8x8_wrap mul_252(.CLK(CLK), .W(W[2023:2016]), .IMG(IMG[2023:2016]), .P(mul_out_252));
   mul8x8_wrap mul_253(.CLK(CLK), .W(W[2031:2024]), .IMG(IMG[2031:2024]), .P(mul_out_253));
   mul8x8_wrap mul_254(.CLK(CLK), .W(W[2039:2032]), .IMG(IMG[2039:2032]), .P(mul_out_254));
   mul8x8_wrap mul_255(.CLK(CLK), .W(W[2047:2040]), .IMG(IMG[2047:2040]), .P(mul_out_255));
   mul8x8_wrap mul_256(.CLK(CLK), .W(W[2055:2048]), .IMG(IMG[2055:2048]), .P(mul_out_256));
   mul8x8_wrap mul_257(.CLK(CLK), .W(W[2063:2056]), .IMG(IMG[2063:2056]), .P(mul_out_257));
   mul8x8_wrap mul_258(.CLK(CLK), .W(W[2071:2064]), .IMG(IMG[2071:2064]), .P(mul_out_258));
   mul8x8_wrap mul_259(.CLK(CLK), .W(W[2079:2072]), .IMG(IMG[2079:2072]), .P(mul_out_259));
   mul8x8_wrap mul_260(.CLK(CLK), .W(W[2087:2080]), .IMG(IMG[2087:2080]), .P(mul_out_260));
   mul8x8_wrap mul_261(.CLK(CLK), .W(W[2095:2088]), .IMG(IMG[2095:2088]), .P(mul_out_261));
   mul8x8_wrap mul_262(.CLK(CLK), .W(W[2103:2096]), .IMG(IMG[2103:2096]), .P(mul_out_262));
   mul8x8_wrap mul_263(.CLK(CLK), .W(W[2111:2104]), .IMG(IMG[2111:2104]), .P(mul_out_263));
   mul8x8_wrap mul_264(.CLK(CLK), .W(W[2119:2112]), .IMG(IMG[2119:2112]), .P(mul_out_264));
   mul8x8_wrap mul_265(.CLK(CLK), .W(W[2127:2120]), .IMG(IMG[2127:2120]), .P(mul_out_265));
   mul8x8_wrap mul_266(.CLK(CLK), .W(W[2135:2128]), .IMG(IMG[2135:2128]), .P(mul_out_266));
   mul8x8_wrap mul_267(.CLK(CLK), .W(W[2143:2136]), .IMG(IMG[2143:2136]), .P(mul_out_267));
   mul8x8_wrap mul_268(.CLK(CLK), .W(W[2151:2144]), .IMG(IMG[2151:2144]), .P(mul_out_268));
   mul8x8_wrap mul_269(.CLK(CLK), .W(W[2159:2152]), .IMG(IMG[2159:2152]), .P(mul_out_269));
   mul8x8_wrap mul_270(.CLK(CLK), .W(W[2167:2160]), .IMG(IMG[2167:2160]), .P(mul_out_270));
   mul8x8_wrap mul_271(.CLK(CLK), .W(W[2175:2168]), .IMG(IMG[2175:2168]), .P(mul_out_271));
   mul8x8_wrap mul_272(.CLK(CLK), .W(W[2183:2176]), .IMG(IMG[2183:2176]), .P(mul_out_272));
   mul8x8_wrap mul_273(.CLK(CLK), .W(W[2191:2184]), .IMG(IMG[2191:2184]), .P(mul_out_273));
   mul8x8_wrap mul_274(.CLK(CLK), .W(W[2199:2192]), .IMG(IMG[2199:2192]), .P(mul_out_274));
   mul8x8_wrap mul_275(.CLK(CLK), .W(W[2207:2200]), .IMG(IMG[2207:2200]), .P(mul_out_275));
   mul8x8_wrap mul_276(.CLK(CLK), .W(W[2215:2208]), .IMG(IMG[2215:2208]), .P(mul_out_276));
   mul8x8_wrap mul_277(.CLK(CLK), .W(W[2223:2216]), .IMG(IMG[2223:2216]), .P(mul_out_277));
   mul8x8_wrap mul_278(.CLK(CLK), .W(W[2231:2224]), .IMG(IMG[2231:2224]), .P(mul_out_278));
   mul8x8_wrap mul_279(.CLK(CLK), .W(W[2239:2232]), .IMG(IMG[2239:2232]), .P(mul_out_279));
   mul8x8_wrap mul_280(.CLK(CLK), .W(W[2247:2240]), .IMG(IMG[2247:2240]), .P(mul_out_280));
   mul8x8_wrap mul_281(.CLK(CLK), .W(W[2255:2248]), .IMG(IMG[2255:2248]), .P(mul_out_281));
   mul8x8_wrap mul_282(.CLK(CLK), .W(W[2263:2256]), .IMG(IMG[2263:2256]), .P(mul_out_282));
   mul8x8_wrap mul_283(.CLK(CLK), .W(W[2271:2264]), .IMG(IMG[2271:2264]), .P(mul_out_283));
   mul8x8_wrap mul_284(.CLK(CLK), .W(W[2279:2272]), .IMG(IMG[2279:2272]), .P(mul_out_284));
   mul8x8_wrap mul_285(.CLK(CLK), .W(W[2287:2280]), .IMG(IMG[2287:2280]), .P(mul_out_285));
   mul8x8_wrap mul_286(.CLK(CLK), .W(W[2295:2288]), .IMG(IMG[2295:2288]), .P(mul_out_286));
   mul8x8_wrap mul_287(.CLK(CLK), .W(W[2303:2296]), .IMG(IMG[2303:2296]), .P(mul_out_287));
   mul8x8_wrap mul_288(.CLK(CLK), .W(W[2311:2304]), .IMG(IMG[2311:2304]), .P(mul_out_288));
   mul8x8_wrap mul_289(.CLK(CLK), .W(W[2319:2312]), .IMG(IMG[2319:2312]), .P(mul_out_289));
   mul8x8_wrap mul_290(.CLK(CLK), .W(W[2327:2320]), .IMG(IMG[2327:2320]), .P(mul_out_290));
   mul8x8_wrap mul_291(.CLK(CLK), .W(W[2335:2328]), .IMG(IMG[2335:2328]), .P(mul_out_291));
   mul8x8_wrap mul_292(.CLK(CLK), .W(W[2343:2336]), .IMG(IMG[2343:2336]), .P(mul_out_292));
   mul8x8_wrap mul_293(.CLK(CLK), .W(W[2351:2344]), .IMG(IMG[2351:2344]), .P(mul_out_293));
   mul8x8_wrap mul_294(.CLK(CLK), .W(W[2359:2352]), .IMG(IMG[2359:2352]), .P(mul_out_294));
   mul8x8_wrap mul_295(.CLK(CLK), .W(W[2367:2360]), .IMG(IMG[2367:2360]), .P(mul_out_295));
   mul8x8_wrap mul_296(.CLK(CLK), .W(W[2375:2368]), .IMG(IMG[2375:2368]), .P(mul_out_296));
   mul8x8_wrap mul_297(.CLK(CLK), .W(W[2383:2376]), .IMG(IMG[2383:2376]), .P(mul_out_297));
   mul8x8_wrap mul_298(.CLK(CLK), .W(W[2391:2384]), .IMG(IMG[2391:2384]), .P(mul_out_298));
   mul8x8_wrap mul_299(.CLK(CLK), .W(W[2399:2392]), .IMG(IMG[2399:2392]), .P(mul_out_299));
   mul8x8_wrap mul_300(.CLK(CLK), .W(W[2407:2400]), .IMG(IMG[2407:2400]), .P(mul_out_300));
   mul8x8_wrap mul_301(.CLK(CLK), .W(W[2415:2408]), .IMG(IMG[2415:2408]), .P(mul_out_301));
   mul8x8_wrap mul_302(.CLK(CLK), .W(W[2423:2416]), .IMG(IMG[2423:2416]), .P(mul_out_302));
   mul8x8_wrap mul_303(.CLK(CLK), .W(W[2431:2424]), .IMG(IMG[2431:2424]), .P(mul_out_303));
   mul8x8_wrap mul_304(.CLK(CLK), .W(W[2439:2432]), .IMG(IMG[2439:2432]), .P(mul_out_304));
   mul8x8_wrap mul_305(.CLK(CLK), .W(W[2447:2440]), .IMG(IMG[2447:2440]), .P(mul_out_305));
   mul8x8_wrap mul_306(.CLK(CLK), .W(W[2455:2448]), .IMG(IMG[2455:2448]), .P(mul_out_306));
   mul8x8_wrap mul_307(.CLK(CLK), .W(W[2463:2456]), .IMG(IMG[2463:2456]), .P(mul_out_307));
   mul8x8_wrap mul_308(.CLK(CLK), .W(W[2471:2464]), .IMG(IMG[2471:2464]), .P(mul_out_308));
   mul8x8_wrap mul_309(.CLK(CLK), .W(W[2479:2472]), .IMG(IMG[2479:2472]), .P(mul_out_309));
   mul8x8_wrap mul_310(.CLK(CLK), .W(W[2487:2480]), .IMG(IMG[2487:2480]), .P(mul_out_310));
   mul8x8_wrap mul_311(.CLK(CLK), .W(W[2495:2488]), .IMG(IMG[2495:2488]), .P(mul_out_311));
   mul8x8_wrap mul_312(.CLK(CLK), .W(W[2503:2496]), .IMG(IMG[2503:2496]), .P(mul_out_312));
   mul8x8_wrap mul_313(.CLK(CLK), .W(W[2511:2504]), .IMG(IMG[2511:2504]), .P(mul_out_313));
   mul8x8_wrap mul_314(.CLK(CLK), .W(W[2519:2512]), .IMG(IMG[2519:2512]), .P(mul_out_314));
   mul8x8_wrap mul_315(.CLK(CLK), .W(W[2527:2520]), .IMG(IMG[2527:2520]), .P(mul_out_315));
   mul8x8_wrap mul_316(.CLK(CLK), .W(W[2535:2528]), .IMG(IMG[2535:2528]), .P(mul_out_316));
   mul8x8_wrap mul_317(.CLK(CLK), .W(W[2543:2536]), .IMG(IMG[2543:2536]), .P(mul_out_317));
   mul8x8_wrap mul_318(.CLK(CLK), .W(W[2551:2544]), .IMG(IMG[2551:2544]), .P(mul_out_318));
   mul8x8_wrap mul_319(.CLK(CLK), .W(W[2559:2552]), .IMG(IMG[2559:2552]), .P(mul_out_319));
   mul8x8_wrap mul_320(.CLK(CLK), .W(W[2567:2560]), .IMG(IMG[2567:2560]), .P(mul_out_320));
   mul8x8_wrap mul_321(.CLK(CLK), .W(W[2575:2568]), .IMG(IMG[2575:2568]), .P(mul_out_321));
   mul8x8_wrap mul_322(.CLK(CLK), .W(W[2583:2576]), .IMG(IMG[2583:2576]), .P(mul_out_322));
   mul8x8_wrap mul_323(.CLK(CLK), .W(W[2591:2584]), .IMG(IMG[2591:2584]), .P(mul_out_323));
   mul8x8_wrap mul_324(.CLK(CLK), .W(W[2599:2592]), .IMG(IMG[2599:2592]), .P(mul_out_324));
   mul8x8_wrap mul_325(.CLK(CLK), .W(W[2607:2600]), .IMG(IMG[2607:2600]), .P(mul_out_325));
   mul8x8_wrap mul_326(.CLK(CLK), .W(W[2615:2608]), .IMG(IMG[2615:2608]), .P(mul_out_326));
   mul8x8_wrap mul_327(.CLK(CLK), .W(W[2623:2616]), .IMG(IMG[2623:2616]), .P(mul_out_327));
   mul8x8_wrap mul_328(.CLK(CLK), .W(W[2631:2624]), .IMG(IMG[2631:2624]), .P(mul_out_328));
   mul8x8_wrap mul_329(.CLK(CLK), .W(W[2639:2632]), .IMG(IMG[2639:2632]), .P(mul_out_329));
   mul8x8_wrap mul_330(.CLK(CLK), .W(W[2647:2640]), .IMG(IMG[2647:2640]), .P(mul_out_330));
   mul8x8_wrap mul_331(.CLK(CLK), .W(W[2655:2648]), .IMG(IMG[2655:2648]), .P(mul_out_331));
   mul8x8_wrap mul_332(.CLK(CLK), .W(W[2663:2656]), .IMG(IMG[2663:2656]), .P(mul_out_332));
   mul8x8_wrap mul_333(.CLK(CLK), .W(W[2671:2664]), .IMG(IMG[2671:2664]), .P(mul_out_333));
   mul8x8_wrap mul_334(.CLK(CLK), .W(W[2679:2672]), .IMG(IMG[2679:2672]), .P(mul_out_334));
   mul8x8_wrap mul_335(.CLK(CLK), .W(W[2687:2680]), .IMG(IMG[2687:2680]), .P(mul_out_335));
   mul8x8_wrap mul_336(.CLK(CLK), .W(W[2695:2688]), .IMG(IMG[2695:2688]), .P(mul_out_336));
   mul8x8_wrap mul_337(.CLK(CLK), .W(W[2703:2696]), .IMG(IMG[2703:2696]), .P(mul_out_337));
   mul8x8_wrap mul_338(.CLK(CLK), .W(W[2711:2704]), .IMG(IMG[2711:2704]), .P(mul_out_338));
   mul8x8_wrap mul_339(.CLK(CLK), .W(W[2719:2712]), .IMG(IMG[2719:2712]), .P(mul_out_339));
   mul8x8_wrap mul_340(.CLK(CLK), .W(W[2727:2720]), .IMG(IMG[2727:2720]), .P(mul_out_340));
   mul8x8_wrap mul_341(.CLK(CLK), .W(W[2735:2728]), .IMG(IMG[2735:2728]), .P(mul_out_341));
   mul8x8_wrap mul_342(.CLK(CLK), .W(W[2743:2736]), .IMG(IMG[2743:2736]), .P(mul_out_342));
   mul8x8_wrap mul_343(.CLK(CLK), .W(W[2751:2744]), .IMG(IMG[2751:2744]), .P(mul_out_343));
   mul8x8_wrap mul_344(.CLK(CLK), .W(W[2759:2752]), .IMG(IMG[2759:2752]), .P(mul_out_344));
   mul8x8_wrap mul_345(.CLK(CLK), .W(W[2767:2760]), .IMG(IMG[2767:2760]), .P(mul_out_345));
   mul8x8_wrap mul_346(.CLK(CLK), .W(W[2775:2768]), .IMG(IMG[2775:2768]), .P(mul_out_346));
   mul8x8_wrap mul_347(.CLK(CLK), .W(W[2783:2776]), .IMG(IMG[2783:2776]), .P(mul_out_347));
   mul8x8_wrap mul_348(.CLK(CLK), .W(W[2791:2784]), .IMG(IMG[2791:2784]), .P(mul_out_348));
   mul8x8_wrap mul_349(.CLK(CLK), .W(W[2799:2792]), .IMG(IMG[2799:2792]), .P(mul_out_349));
   mul8x8_wrap mul_350(.CLK(CLK), .W(W[2807:2800]), .IMG(IMG[2807:2800]), .P(mul_out_350));
   mul8x8_wrap mul_351(.CLK(CLK), .W(W[2815:2808]), .IMG(IMG[2815:2808]), .P(mul_out_351));
   mul8x8_wrap mul_352(.CLK(CLK), .W(W[2823:2816]), .IMG(IMG[2823:2816]), .P(mul_out_352));
   mul8x8_wrap mul_353(.CLK(CLK), .W(W[2831:2824]), .IMG(IMG[2831:2824]), .P(mul_out_353));
   mul8x8_wrap mul_354(.CLK(CLK), .W(W[2839:2832]), .IMG(IMG[2839:2832]), .P(mul_out_354));
   mul8x8_wrap mul_355(.CLK(CLK), .W(W[2847:2840]), .IMG(IMG[2847:2840]), .P(mul_out_355));
   mul8x8_wrap mul_356(.CLK(CLK), .W(W[2855:2848]), .IMG(IMG[2855:2848]), .P(mul_out_356));
   mul8x8_wrap mul_357(.CLK(CLK), .W(W[2863:2856]), .IMG(IMG[2863:2856]), .P(mul_out_357));
   mul8x8_wrap mul_358(.CLK(CLK), .W(W[2871:2864]), .IMG(IMG[2871:2864]), .P(mul_out_358));
   mul8x8_wrap mul_359(.CLK(CLK), .W(W[2879:2872]), .IMG(IMG[2879:2872]), .P(mul_out_359));
   mul8x8_wrap mul_360(.CLK(CLK), .W(W[2887:2880]), .IMG(IMG[2887:2880]), .P(mul_out_360));
   mul8x8_wrap mul_361(.CLK(CLK), .W(W[2895:2888]), .IMG(IMG[2895:2888]), .P(mul_out_361));
   mul8x8_wrap mul_362(.CLK(CLK), .W(W[2903:2896]), .IMG(IMG[2903:2896]), .P(mul_out_362));
   mul8x8_wrap mul_363(.CLK(CLK), .W(W[2911:2904]), .IMG(IMG[2911:2904]), .P(mul_out_363));
   mul8x8_wrap mul_364(.CLK(CLK), .W(W[2919:2912]), .IMG(IMG[2919:2912]), .P(mul_out_364));
   mul8x8_wrap mul_365(.CLK(CLK), .W(W[2927:2920]), .IMG(IMG[2927:2920]), .P(mul_out_365));
   mul8x8_wrap mul_366(.CLK(CLK), .W(W[2935:2928]), .IMG(IMG[2935:2928]), .P(mul_out_366));
   mul8x8_wrap mul_367(.CLK(CLK), .W(W[2943:2936]), .IMG(IMG[2943:2936]), .P(mul_out_367));
   mul8x8_wrap mul_368(.CLK(CLK), .W(W[2951:2944]), .IMG(IMG[2951:2944]), .P(mul_out_368));
   mul8x8_wrap mul_369(.CLK(CLK), .W(W[2959:2952]), .IMG(IMG[2959:2952]), .P(mul_out_369));
   mul8x8_wrap mul_370(.CLK(CLK), .W(W[2967:2960]), .IMG(IMG[2967:2960]), .P(mul_out_370));
   mul8x8_wrap mul_371(.CLK(CLK), .W(W[2975:2968]), .IMG(IMG[2975:2968]), .P(mul_out_371));
   mul8x8_wrap mul_372(.CLK(CLK), .W(W[2983:2976]), .IMG(IMG[2983:2976]), .P(mul_out_372));
   mul8x8_wrap mul_373(.CLK(CLK), .W(W[2991:2984]), .IMG(IMG[2991:2984]), .P(mul_out_373));
   mul8x8_wrap mul_374(.CLK(CLK), .W(W[2999:2992]), .IMG(IMG[2999:2992]), .P(mul_out_374));
   mul8x8_wrap mul_375(.CLK(CLK), .W(W[3007:3000]), .IMG(IMG[3007:3000]), .P(mul_out_375));
   mul8x8_wrap mul_376(.CLK(CLK), .W(W[3015:3008]), .IMG(IMG[3015:3008]), .P(mul_out_376));
   mul8x8_wrap mul_377(.CLK(CLK), .W(W[3023:3016]), .IMG(IMG[3023:3016]), .P(mul_out_377));
   mul8x8_wrap mul_378(.CLK(CLK), .W(W[3031:3024]), .IMG(IMG[3031:3024]), .P(mul_out_378));
   mul8x8_wrap mul_379(.CLK(CLK), .W(W[3039:3032]), .IMG(IMG[3039:3032]), .P(mul_out_379));
   mul8x8_wrap mul_380(.CLK(CLK), .W(W[3047:3040]), .IMG(IMG[3047:3040]), .P(mul_out_380));
   mul8x8_wrap mul_381(.CLK(CLK), .W(W[3055:3048]), .IMG(IMG[3055:3048]), .P(mul_out_381));
   mul8x8_wrap mul_382(.CLK(CLK), .W(W[3063:3056]), .IMG(IMG[3063:3056]), .P(mul_out_382));
   mul8x8_wrap mul_383(.CLK(CLK), .W(W[3071:3064]), .IMG(IMG[3071:3064]), .P(mul_out_383));
   mul8x8_wrap mul_384(.CLK(CLK), .W(W[3079:3072]), .IMG(IMG[3079:3072]), .P(mul_out_384));
   mul8x8_wrap mul_385(.CLK(CLK), .W(W[3087:3080]), .IMG(IMG[3087:3080]), .P(mul_out_385));
   mul8x8_wrap mul_386(.CLK(CLK), .W(W[3095:3088]), .IMG(IMG[3095:3088]), .P(mul_out_386));
   mul8x8_wrap mul_387(.CLK(CLK), .W(W[3103:3096]), .IMG(IMG[3103:3096]), .P(mul_out_387));
   mul8x8_wrap mul_388(.CLK(CLK), .W(W[3111:3104]), .IMG(IMG[3111:3104]), .P(mul_out_388));
   mul8x8_wrap mul_389(.CLK(CLK), .W(W[3119:3112]), .IMG(IMG[3119:3112]), .P(mul_out_389));
   mul8x8_wrap mul_390(.CLK(CLK), .W(W[3127:3120]), .IMG(IMG[3127:3120]), .P(mul_out_390));
   mul8x8_wrap mul_391(.CLK(CLK), .W(W[3135:3128]), .IMG(IMG[3135:3128]), .P(mul_out_391));
   mul8x8_wrap mul_392(.CLK(CLK), .W(W[3143:3136]), .IMG(IMG[3143:3136]), .P(mul_out_392));
   mul8x8_wrap mul_393(.CLK(CLK), .W(W[3151:3144]), .IMG(IMG[3151:3144]), .P(mul_out_393));
   mul8x8_wrap mul_394(.CLK(CLK), .W(W[3159:3152]), .IMG(IMG[3159:3152]), .P(mul_out_394));
   mul8x8_wrap mul_395(.CLK(CLK), .W(W[3167:3160]), .IMG(IMG[3167:3160]), .P(mul_out_395));
   mul8x8_wrap mul_396(.CLK(CLK), .W(W[3175:3168]), .IMG(IMG[3175:3168]), .P(mul_out_396));
   mul8x8_wrap mul_397(.CLK(CLK), .W(W[3183:3176]), .IMG(IMG[3183:3176]), .P(mul_out_397));
   mul8x8_wrap mul_398(.CLK(CLK), .W(W[3191:3184]), .IMG(IMG[3191:3184]), .P(mul_out_398));
   mul8x8_wrap mul_399(.CLK(CLK), .W(W[3199:3192]), .IMG(IMG[3199:3192]), .P(mul_out_399));
   mul8x8_wrap mul_400(.CLK(CLK), .W(W[3207:3200]), .IMG(IMG[3207:3200]), .P(mul_out_400));
   mul8x8_wrap mul_401(.CLK(CLK), .W(W[3215:3208]), .IMG(IMG[3215:3208]), .P(mul_out_401));
   mul8x8_wrap mul_402(.CLK(CLK), .W(W[3223:3216]), .IMG(IMG[3223:3216]), .P(mul_out_402));
   mul8x8_wrap mul_403(.CLK(CLK), .W(W[3231:3224]), .IMG(IMG[3231:3224]), .P(mul_out_403));
   mul8x8_wrap mul_404(.CLK(CLK), .W(W[3239:3232]), .IMG(IMG[3239:3232]), .P(mul_out_404));
   mul8x8_wrap mul_405(.CLK(CLK), .W(W[3247:3240]), .IMG(IMG[3247:3240]), .P(mul_out_405));
   mul8x8_wrap mul_406(.CLK(CLK), .W(W[3255:3248]), .IMG(IMG[3255:3248]), .P(mul_out_406));
   mul8x8_wrap mul_407(.CLK(CLK), .W(W[3263:3256]), .IMG(IMG[3263:3256]), .P(mul_out_407));
   mul8x8_wrap mul_408(.CLK(CLK), .W(W[3271:3264]), .IMG(IMG[3271:3264]), .P(mul_out_408));
   mul8x8_wrap mul_409(.CLK(CLK), .W(W[3279:3272]), .IMG(IMG[3279:3272]), .P(mul_out_409));
   mul8x8_wrap mul_410(.CLK(CLK), .W(W[3287:3280]), .IMG(IMG[3287:3280]), .P(mul_out_410));
   mul8x8_wrap mul_411(.CLK(CLK), .W(W[3295:3288]), .IMG(IMG[3295:3288]), .P(mul_out_411));
   mul8x8_wrap mul_412(.CLK(CLK), .W(W[3303:3296]), .IMG(IMG[3303:3296]), .P(mul_out_412));
   mul8x8_wrap mul_413(.CLK(CLK), .W(W[3311:3304]), .IMG(IMG[3311:3304]), .P(mul_out_413));
   mul8x8_wrap mul_414(.CLK(CLK), .W(W[3319:3312]), .IMG(IMG[3319:3312]), .P(mul_out_414));
   mul8x8_wrap mul_415(.CLK(CLK), .W(W[3327:3320]), .IMG(IMG[3327:3320]), .P(mul_out_415));
   mul8x8_wrap mul_416(.CLK(CLK), .W(W[3335:3328]), .IMG(IMG[3335:3328]), .P(mul_out_416));
   mul8x8_wrap mul_417(.CLK(CLK), .W(W[3343:3336]), .IMG(IMG[3343:3336]), .P(mul_out_417));
   mul8x8_wrap mul_418(.CLK(CLK), .W(W[3351:3344]), .IMG(IMG[3351:3344]), .P(mul_out_418));
   mul8x8_wrap mul_419(.CLK(CLK), .W(W[3359:3352]), .IMG(IMG[3359:3352]), .P(mul_out_419));
   mul8x8_wrap mul_420(.CLK(CLK), .W(W[3367:3360]), .IMG(IMG[3367:3360]), .P(mul_out_420));
   mul8x8_wrap mul_421(.CLK(CLK), .W(W[3375:3368]), .IMG(IMG[3375:3368]), .P(mul_out_421));
   mul8x8_wrap mul_422(.CLK(CLK), .W(W[3383:3376]), .IMG(IMG[3383:3376]), .P(mul_out_422));
   mul8x8_wrap mul_423(.CLK(CLK), .W(W[3391:3384]), .IMG(IMG[3391:3384]), .P(mul_out_423));
   mul8x8_wrap mul_424(.CLK(CLK), .W(W[3399:3392]), .IMG(IMG[3399:3392]), .P(mul_out_424));
   mul8x8_wrap mul_425(.CLK(CLK), .W(W[3407:3400]), .IMG(IMG[3407:3400]), .P(mul_out_425));
   mul8x8_wrap mul_426(.CLK(CLK), .W(W[3415:3408]), .IMG(IMG[3415:3408]), .P(mul_out_426));
   mul8x8_wrap mul_427(.CLK(CLK), .W(W[3423:3416]), .IMG(IMG[3423:3416]), .P(mul_out_427));
   mul8x8_wrap mul_428(.CLK(CLK), .W(W[3431:3424]), .IMG(IMG[3431:3424]), .P(mul_out_428));
   mul8x8_wrap mul_429(.CLK(CLK), .W(W[3439:3432]), .IMG(IMG[3439:3432]), .P(mul_out_429));
   mul8x8_wrap mul_430(.CLK(CLK), .W(W[3447:3440]), .IMG(IMG[3447:3440]), .P(mul_out_430));
   mul8x8_wrap mul_431(.CLK(CLK), .W(W[3455:3448]), .IMG(IMG[3455:3448]), .P(mul_out_431));
   mul8x8_wrap mul_432(.CLK(CLK), .W(W[3463:3456]), .IMG(IMG[3463:3456]), .P(mul_out_432));
   mul8x8_wrap mul_433(.CLK(CLK), .W(W[3471:3464]), .IMG(IMG[3471:3464]), .P(mul_out_433));
   mul8x8_wrap mul_434(.CLK(CLK), .W(W[3479:3472]), .IMG(IMG[3479:3472]), .P(mul_out_434));
   mul8x8_wrap mul_435(.CLK(CLK), .W(W[3487:3480]), .IMG(IMG[3487:3480]), .P(mul_out_435));
   mul8x8_wrap mul_436(.CLK(CLK), .W(W[3495:3488]), .IMG(IMG[3495:3488]), .P(mul_out_436));
   mul8x8_wrap mul_437(.CLK(CLK), .W(W[3503:3496]), .IMG(IMG[3503:3496]), .P(mul_out_437));
   mul8x8_wrap mul_438(.CLK(CLK), .W(W[3511:3504]), .IMG(IMG[3511:3504]), .P(mul_out_438));
   mul8x8_wrap mul_439(.CLK(CLK), .W(W[3519:3512]), .IMG(IMG[3519:3512]), .P(mul_out_439));
   mul8x8_wrap mul_440(.CLK(CLK), .W(W[3527:3520]), .IMG(IMG[3527:3520]), .P(mul_out_440));
   mul8x8_wrap mul_441(.CLK(CLK), .W(W[3535:3528]), .IMG(IMG[3535:3528]), .P(mul_out_441));
   mul8x8_wrap mul_442(.CLK(CLK), .W(W[3543:3536]), .IMG(IMG[3543:3536]), .P(mul_out_442));
   mul8x8_wrap mul_443(.CLK(CLK), .W(W[3551:3544]), .IMG(IMG[3551:3544]), .P(mul_out_443));
   mul8x8_wrap mul_444(.CLK(CLK), .W(W[3559:3552]), .IMG(IMG[3559:3552]), .P(mul_out_444));
   mul8x8_wrap mul_445(.CLK(CLK), .W(W[3567:3560]), .IMG(IMG[3567:3560]), .P(mul_out_445));
   mul8x8_wrap mul_446(.CLK(CLK), .W(W[3575:3568]), .IMG(IMG[3575:3568]), .P(mul_out_446));
   mul8x8_wrap mul_447(.CLK(CLK), .W(W[3583:3576]), .IMG(IMG[3583:3576]), .P(mul_out_447));
   mul8x8_wrap mul_448(.CLK(CLK), .W(W[3591:3584]), .IMG(IMG[3591:3584]), .P(mul_out_448));
   mul8x8_wrap mul_449(.CLK(CLK), .W(W[3599:3592]), .IMG(IMG[3599:3592]), .P(mul_out_449));
   mul8x8_wrap mul_450(.CLK(CLK), .W(W[3607:3600]), .IMG(IMG[3607:3600]), .P(mul_out_450));
   mul8x8_wrap mul_451(.CLK(CLK), .W(W[3615:3608]), .IMG(IMG[3615:3608]), .P(mul_out_451));
   mul8x8_wrap mul_452(.CLK(CLK), .W(W[3623:3616]), .IMG(IMG[3623:3616]), .P(mul_out_452));
   mul8x8_wrap mul_453(.CLK(CLK), .W(W[3631:3624]), .IMG(IMG[3631:3624]), .P(mul_out_453));
   mul8x8_wrap mul_454(.CLK(CLK), .W(W[3639:3632]), .IMG(IMG[3639:3632]), .P(mul_out_454));
   mul8x8_wrap mul_455(.CLK(CLK), .W(W[3647:3640]), .IMG(IMG[3647:3640]), .P(mul_out_455));
   mul8x8_wrap mul_456(.CLK(CLK), .W(W[3655:3648]), .IMG(IMG[3655:3648]), .P(mul_out_456));
   mul8x8_wrap mul_457(.CLK(CLK), .W(W[3663:3656]), .IMG(IMG[3663:3656]), .P(mul_out_457));
   mul8x8_wrap mul_458(.CLK(CLK), .W(W[3671:3664]), .IMG(IMG[3671:3664]), .P(mul_out_458));
   mul8x8_wrap mul_459(.CLK(CLK), .W(W[3679:3672]), .IMG(IMG[3679:3672]), .P(mul_out_459));
   mul8x8_wrap mul_460(.CLK(CLK), .W(W[3687:3680]), .IMG(IMG[3687:3680]), .P(mul_out_460));
   mul8x8_wrap mul_461(.CLK(CLK), .W(W[3695:3688]), .IMG(IMG[3695:3688]), .P(mul_out_461));
   mul8x8_wrap mul_462(.CLK(CLK), .W(W[3703:3696]), .IMG(IMG[3703:3696]), .P(mul_out_462));
   mul8x8_wrap mul_463(.CLK(CLK), .W(W[3711:3704]), .IMG(IMG[3711:3704]), .P(mul_out_463));
   mul8x8_wrap mul_464(.CLK(CLK), .W(W[3719:3712]), .IMG(IMG[3719:3712]), .P(mul_out_464));
   mul8x8_wrap mul_465(.CLK(CLK), .W(W[3727:3720]), .IMG(IMG[3727:3720]), .P(mul_out_465));
   mul8x8_wrap mul_466(.CLK(CLK), .W(W[3735:3728]), .IMG(IMG[3735:3728]), .P(mul_out_466));
   mul8x8_wrap mul_467(.CLK(CLK), .W(W[3743:3736]), .IMG(IMG[3743:3736]), .P(mul_out_467));
   mul8x8_wrap mul_468(.CLK(CLK), .W(W[3751:3744]), .IMG(IMG[3751:3744]), .P(mul_out_468));
   mul8x8_wrap mul_469(.CLK(CLK), .W(W[3759:3752]), .IMG(IMG[3759:3752]), .P(mul_out_469));
   mul8x8_wrap mul_470(.CLK(CLK), .W(W[3767:3760]), .IMG(IMG[3767:3760]), .P(mul_out_470));
   mul8x8_wrap mul_471(.CLK(CLK), .W(W[3775:3768]), .IMG(IMG[3775:3768]), .P(mul_out_471));
   mul8x8_wrap mul_472(.CLK(CLK), .W(W[3783:3776]), .IMG(IMG[3783:3776]), .P(mul_out_472));
   mul8x8_wrap mul_473(.CLK(CLK), .W(W[3791:3784]), .IMG(IMG[3791:3784]), .P(mul_out_473));
   mul8x8_wrap mul_474(.CLK(CLK), .W(W[3799:3792]), .IMG(IMG[3799:3792]), .P(mul_out_474));
   mul8x8_wrap mul_475(.CLK(CLK), .W(W[3807:3800]), .IMG(IMG[3807:3800]), .P(mul_out_475));
   mul8x8_wrap mul_476(.CLK(CLK), .W(W[3815:3808]), .IMG(IMG[3815:3808]), .P(mul_out_476));
   mul8x8_wrap mul_477(.CLK(CLK), .W(W[3823:3816]), .IMG(IMG[3823:3816]), .P(mul_out_477));
   mul8x8_wrap mul_478(.CLK(CLK), .W(W[3831:3824]), .IMG(IMG[3831:3824]), .P(mul_out_478));
   mul8x8_wrap mul_479(.CLK(CLK), .W(W[3839:3832]), .IMG(IMG[3839:3832]), .P(mul_out_479));
   mul8x8_wrap mul_480(.CLK(CLK), .W(W[3847:3840]), .IMG(IMG[3847:3840]), .P(mul_out_480));
   mul8x8_wrap mul_481(.CLK(CLK), .W(W[3855:3848]), .IMG(IMG[3855:3848]), .P(mul_out_481));
   mul8x8_wrap mul_482(.CLK(CLK), .W(W[3863:3856]), .IMG(IMG[3863:3856]), .P(mul_out_482));
   mul8x8_wrap mul_483(.CLK(CLK), .W(W[3871:3864]), .IMG(IMG[3871:3864]), .P(mul_out_483));
   mul8x8_wrap mul_484(.CLK(CLK), .W(W[3879:3872]), .IMG(IMG[3879:3872]), .P(mul_out_484));
   mul8x8_wrap mul_485(.CLK(CLK), .W(W[3887:3880]), .IMG(IMG[3887:3880]), .P(mul_out_485));
   mul8x8_wrap mul_486(.CLK(CLK), .W(W[3895:3888]), .IMG(IMG[3895:3888]), .P(mul_out_486));
   mul8x8_wrap mul_487(.CLK(CLK), .W(W[3903:3896]), .IMG(IMG[3903:3896]), .P(mul_out_487));
   mul8x8_wrap mul_488(.CLK(CLK), .W(W[3911:3904]), .IMG(IMG[3911:3904]), .P(mul_out_488));
   mul8x8_wrap mul_489(.CLK(CLK), .W(W[3919:3912]), .IMG(IMG[3919:3912]), .P(mul_out_489));
   mul8x8_wrap mul_490(.CLK(CLK), .W(W[3927:3920]), .IMG(IMG[3927:3920]), .P(mul_out_490));
   mul8x8_wrap mul_491(.CLK(CLK), .W(W[3935:3928]), .IMG(IMG[3935:3928]), .P(mul_out_491));
   mul8x8_wrap mul_492(.CLK(CLK), .W(W[3943:3936]), .IMG(IMG[3943:3936]), .P(mul_out_492));
   mul8x8_wrap mul_493(.CLK(CLK), .W(W[3951:3944]), .IMG(IMG[3951:3944]), .P(mul_out_493));
   mul8x8_wrap mul_494(.CLK(CLK), .W(W[3959:3952]), .IMG(IMG[3959:3952]), .P(mul_out_494));
   mul8x8_wrap mul_495(.CLK(CLK), .W(W[3967:3960]), .IMG(IMG[3967:3960]), .P(mul_out_495));
   mul8x8_wrap mul_496(.CLK(CLK), .W(W[3975:3968]), .IMG(IMG[3975:3968]), .P(mul_out_496));
   mul8x8_wrap mul_497(.CLK(CLK), .W(W[3983:3976]), .IMG(IMG[3983:3976]), .P(mul_out_497));
   mul8x8_wrap mul_498(.CLK(CLK), .W(W[3991:3984]), .IMG(IMG[3991:3984]), .P(mul_out_498));
   mul8x8_wrap mul_499(.CLK(CLK), .W(W[3999:3992]), .IMG(IMG[3999:3992]), .P(mul_out_499));
   mul8x8_wrap mul_500(.CLK(CLK), .W(W[4007:4000]), .IMG(IMG[4007:4000]), .P(mul_out_500));
   mul8x8_wrap mul_501(.CLK(CLK), .W(W[4015:4008]), .IMG(IMG[4015:4008]), .P(mul_out_501));
   mul8x8_wrap mul_502(.CLK(CLK), .W(W[4023:4016]), .IMG(IMG[4023:4016]), .P(mul_out_502));
   mul8x8_wrap mul_503(.CLK(CLK), .W(W[4031:4024]), .IMG(IMG[4031:4024]), .P(mul_out_503));
   mul8x8_wrap mul_504(.CLK(CLK), .W(W[4039:4032]), .IMG(IMG[4039:4032]), .P(mul_out_504));
   mul8x8_wrap mul_505(.CLK(CLK), .W(W[4047:4040]), .IMG(IMG[4047:4040]), .P(mul_out_505));
   mul8x8_wrap mul_506(.CLK(CLK), .W(W[4055:4048]), .IMG(IMG[4055:4048]), .P(mul_out_506));
   mul8x8_wrap mul_507(.CLK(CLK), .W(W[4063:4056]), .IMG(IMG[4063:4056]), .P(mul_out_507));
   mul8x8_wrap mul_508(.CLK(CLK), .W(W[4071:4064]), .IMG(IMG[4071:4064]), .P(mul_out_508));
   mul8x8_wrap mul_509(.CLK(CLK), .W(W[4079:4072]), .IMG(IMG[4079:4072]), .P(mul_out_509));
   mul8x8_wrap mul_510(.CLK(CLK), .W(W[4087:4080]), .IMG(IMG[4087:4080]), .P(mul_out_510));
   mul8x8_wrap mul_511(.CLK(CLK), .W(W[4095:4088]), .IMG(IMG[4095:4088]), .P(mul_out_511));
   mul8x8_wrap mul_512(.CLK(CLK), .W(W[4103:4096]), .IMG(IMG[4103:4096]), .P(mul_out_512));
   mul8x8_wrap mul_513(.CLK(CLK), .W(W[4111:4104]), .IMG(IMG[4111:4104]), .P(mul_out_513));
   mul8x8_wrap mul_514(.CLK(CLK), .W(W[4119:4112]), .IMG(IMG[4119:4112]), .P(mul_out_514));
   mul8x8_wrap mul_515(.CLK(CLK), .W(W[4127:4120]), .IMG(IMG[4127:4120]), .P(mul_out_515));
   mul8x8_wrap mul_516(.CLK(CLK), .W(W[4135:4128]), .IMG(IMG[4135:4128]), .P(mul_out_516));
   mul8x8_wrap mul_517(.CLK(CLK), .W(W[4143:4136]), .IMG(IMG[4143:4136]), .P(mul_out_517));
   mul8x8_wrap mul_518(.CLK(CLK), .W(W[4151:4144]), .IMG(IMG[4151:4144]), .P(mul_out_518));
   mul8x8_wrap mul_519(.CLK(CLK), .W(W[4159:4152]), .IMG(IMG[4159:4152]), .P(mul_out_519));
   mul8x8_wrap mul_520(.CLK(CLK), .W(W[4167:4160]), .IMG(IMG[4167:4160]), .P(mul_out_520));
   mul8x8_wrap mul_521(.CLK(CLK), .W(W[4175:4168]), .IMG(IMG[4175:4168]), .P(mul_out_521));
   mul8x8_wrap mul_522(.CLK(CLK), .W(W[4183:4176]), .IMG(IMG[4183:4176]), .P(mul_out_522));
   mul8x8_wrap mul_523(.CLK(CLK), .W(W[4191:4184]), .IMG(IMG[4191:4184]), .P(mul_out_523));
   mul8x8_wrap mul_524(.CLK(CLK), .W(W[4199:4192]), .IMG(IMG[4199:4192]), .P(mul_out_524));
   mul8x8_wrap mul_525(.CLK(CLK), .W(W[4207:4200]), .IMG(IMG[4207:4200]), .P(mul_out_525));
   mul8x8_wrap mul_526(.CLK(CLK), .W(W[4215:4208]), .IMG(IMG[4215:4208]), .P(mul_out_526));
   mul8x8_wrap mul_527(.CLK(CLK), .W(W[4223:4216]), .IMG(IMG[4223:4216]), .P(mul_out_527));
   mul8x8_wrap mul_528(.CLK(CLK), .W(W[4231:4224]), .IMG(IMG[4231:4224]), .P(mul_out_528));
   mul8x8_wrap mul_529(.CLK(CLK), .W(W[4239:4232]), .IMG(IMG[4239:4232]), .P(mul_out_529));
   mul8x8_wrap mul_530(.CLK(CLK), .W(W[4247:4240]), .IMG(IMG[4247:4240]), .P(mul_out_530));
   mul8x8_wrap mul_531(.CLK(CLK), .W(W[4255:4248]), .IMG(IMG[4255:4248]), .P(mul_out_531));
   mul8x8_wrap mul_532(.CLK(CLK), .W(W[4263:4256]), .IMG(IMG[4263:4256]), .P(mul_out_532));
   mul8x8_wrap mul_533(.CLK(CLK), .W(W[4271:4264]), .IMG(IMG[4271:4264]), .P(mul_out_533));
   mul8x8_wrap mul_534(.CLK(CLK), .W(W[4279:4272]), .IMG(IMG[4279:4272]), .P(mul_out_534));
   mul8x8_wrap mul_535(.CLK(CLK), .W(W[4287:4280]), .IMG(IMG[4287:4280]), .P(mul_out_535));
   mul8x8_wrap mul_536(.CLK(CLK), .W(W[4295:4288]), .IMG(IMG[4295:4288]), .P(mul_out_536));
   mul8x8_wrap mul_537(.CLK(CLK), .W(W[4303:4296]), .IMG(IMG[4303:4296]), .P(mul_out_537));
   mul8x8_wrap mul_538(.CLK(CLK), .W(W[4311:4304]), .IMG(IMG[4311:4304]), .P(mul_out_538));
   mul8x8_wrap mul_539(.CLK(CLK), .W(W[4319:4312]), .IMG(IMG[4319:4312]), .P(mul_out_539));
   mul8x8_wrap mul_540(.CLK(CLK), .W(W[4327:4320]), .IMG(IMG[4327:4320]), .P(mul_out_540));
   mul8x8_wrap mul_541(.CLK(CLK), .W(W[4335:4328]), .IMG(IMG[4335:4328]), .P(mul_out_541));
   mul8x8_wrap mul_542(.CLK(CLK), .W(W[4343:4336]), .IMG(IMG[4343:4336]), .P(mul_out_542));
   mul8x8_wrap mul_543(.CLK(CLK), .W(W[4351:4344]), .IMG(IMG[4351:4344]), .P(mul_out_543));
   mul8x8_wrap mul_544(.CLK(CLK), .W(W[4359:4352]), .IMG(IMG[4359:4352]), .P(mul_out_544));
   mul8x8_wrap mul_545(.CLK(CLK), .W(W[4367:4360]), .IMG(IMG[4367:4360]), .P(mul_out_545));
   mul8x8_wrap mul_546(.CLK(CLK), .W(W[4375:4368]), .IMG(IMG[4375:4368]), .P(mul_out_546));
   mul8x8_wrap mul_547(.CLK(CLK), .W(W[4383:4376]), .IMG(IMG[4383:4376]), .P(mul_out_547));
   mul8x8_wrap mul_548(.CLK(CLK), .W(W[4391:4384]), .IMG(IMG[4391:4384]), .P(mul_out_548));
   mul8x8_wrap mul_549(.CLK(CLK), .W(W[4399:4392]), .IMG(IMG[4399:4392]), .P(mul_out_549));
   mul8x8_wrap mul_550(.CLK(CLK), .W(W[4407:4400]), .IMG(IMG[4407:4400]), .P(mul_out_550));
   mul8x8_wrap mul_551(.CLK(CLK), .W(W[4415:4408]), .IMG(IMG[4415:4408]), .P(mul_out_551));
   mul8x8_wrap mul_552(.CLK(CLK), .W(W[4423:4416]), .IMG(IMG[4423:4416]), .P(mul_out_552));
   mul8x8_wrap mul_553(.CLK(CLK), .W(W[4431:4424]), .IMG(IMG[4431:4424]), .P(mul_out_553));
   mul8x8_wrap mul_554(.CLK(CLK), .W(W[4439:4432]), .IMG(IMG[4439:4432]), .P(mul_out_554));
   mul8x8_wrap mul_555(.CLK(CLK), .W(W[4447:4440]), .IMG(IMG[4447:4440]), .P(mul_out_555));
   mul8x8_wrap mul_556(.CLK(CLK), .W(W[4455:4448]), .IMG(IMG[4455:4448]), .P(mul_out_556));
   mul8x8_wrap mul_557(.CLK(CLK), .W(W[4463:4456]), .IMG(IMG[4463:4456]), .P(mul_out_557));
   mul8x8_wrap mul_558(.CLK(CLK), .W(W[4471:4464]), .IMG(IMG[4471:4464]), .P(mul_out_558));
   mul8x8_wrap mul_559(.CLK(CLK), .W(W[4479:4472]), .IMG(IMG[4479:4472]), .P(mul_out_559));
   mul8x8_wrap mul_560(.CLK(CLK), .W(W[4487:4480]), .IMG(IMG[4487:4480]), .P(mul_out_560));
   mul8x8_wrap mul_561(.CLK(CLK), .W(W[4495:4488]), .IMG(IMG[4495:4488]), .P(mul_out_561));
   mul8x8_wrap mul_562(.CLK(CLK), .W(W[4503:4496]), .IMG(IMG[4503:4496]), .P(mul_out_562));
   mul8x8_wrap mul_563(.CLK(CLK), .W(W[4511:4504]), .IMG(IMG[4511:4504]), .P(mul_out_563));
   mul8x8_wrap mul_564(.CLK(CLK), .W(W[4519:4512]), .IMG(IMG[4519:4512]), .P(mul_out_564));
   mul8x8_wrap mul_565(.CLK(CLK), .W(W[4527:4520]), .IMG(IMG[4527:4520]), .P(mul_out_565));
   mul8x8_wrap mul_566(.CLK(CLK), .W(W[4535:4528]), .IMG(IMG[4535:4528]), .P(mul_out_566));
   mul8x8_wrap mul_567(.CLK(CLK), .W(W[4543:4536]), .IMG(IMG[4543:4536]), .P(mul_out_567));
   mul8x8_wrap mul_568(.CLK(CLK), .W(W[4551:4544]), .IMG(IMG[4551:4544]), .P(mul_out_568));
   mul8x8_wrap mul_569(.CLK(CLK), .W(W[4559:4552]), .IMG(IMG[4559:4552]), .P(mul_out_569));
   mul8x8_wrap mul_570(.CLK(CLK), .W(W[4567:4560]), .IMG(IMG[4567:4560]), .P(mul_out_570));
   mul8x8_wrap mul_571(.CLK(CLK), .W(W[4575:4568]), .IMG(IMG[4575:4568]), .P(mul_out_571));
   mul8x8_wrap mul_572(.CLK(CLK), .W(W[4583:4576]), .IMG(IMG[4583:4576]), .P(mul_out_572));
   mul8x8_wrap mul_573(.CLK(CLK), .W(W[4591:4584]), .IMG(IMG[4591:4584]), .P(mul_out_573));
   mul8x8_wrap mul_574(.CLK(CLK), .W(W[4599:4592]), .IMG(IMG[4599:4592]), .P(mul_out_574));
   mul8x8_wrap mul_575(.CLK(CLK), .W(W[4607:4600]), .IMG(IMG[4607:4600]), .P(mul_out_575));
   mul8x8_wrap mul_576(.CLK(CLK), .W(W[4615:4608]), .IMG(IMG[4615:4608]), .P(mul_out_576));
   mul8x8_wrap mul_577(.CLK(CLK), .W(W[4623:4616]), .IMG(IMG[4623:4616]), .P(mul_out_577));
   mul8x8_wrap mul_578(.CLK(CLK), .W(W[4631:4624]), .IMG(IMG[4631:4624]), .P(mul_out_578));
   mul8x8_wrap mul_579(.CLK(CLK), .W(W[4639:4632]), .IMG(IMG[4639:4632]), .P(mul_out_579));
   mul8x8_wrap mul_580(.CLK(CLK), .W(W[4647:4640]), .IMG(IMG[4647:4640]), .P(mul_out_580));
   mul8x8_wrap mul_581(.CLK(CLK), .W(W[4655:4648]), .IMG(IMG[4655:4648]), .P(mul_out_581));
   mul8x8_wrap mul_582(.CLK(CLK), .W(W[4663:4656]), .IMG(IMG[4663:4656]), .P(mul_out_582));
   mul8x8_wrap mul_583(.CLK(CLK), .W(W[4671:4664]), .IMG(IMG[4671:4664]), .P(mul_out_583));
   mul8x8_wrap mul_584(.CLK(CLK), .W(W[4679:4672]), .IMG(IMG[4679:4672]), .P(mul_out_584));
   mul8x8_wrap mul_585(.CLK(CLK), .W(W[4687:4680]), .IMG(IMG[4687:4680]), .P(mul_out_585));
   mul8x8_wrap mul_586(.CLK(CLK), .W(W[4695:4688]), .IMG(IMG[4695:4688]), .P(mul_out_586));
   mul8x8_wrap mul_587(.CLK(CLK), .W(W[4703:4696]), .IMG(IMG[4703:4696]), .P(mul_out_587));
   mul8x8_wrap mul_588(.CLK(CLK), .W(W[4711:4704]), .IMG(IMG[4711:4704]), .P(mul_out_588));
   mul8x8_wrap mul_589(.CLK(CLK), .W(W[4719:4712]), .IMG(IMG[4719:4712]), .P(mul_out_589));
   mul8x8_wrap mul_590(.CLK(CLK), .W(W[4727:4720]), .IMG(IMG[4727:4720]), .P(mul_out_590));
   mul8x8_wrap mul_591(.CLK(CLK), .W(W[4735:4728]), .IMG(IMG[4735:4728]), .P(mul_out_591));
   mul8x8_wrap mul_592(.CLK(CLK), .W(W[4743:4736]), .IMG(IMG[4743:4736]), .P(mul_out_592));
   mul8x8_wrap mul_593(.CLK(CLK), .W(W[4751:4744]), .IMG(IMG[4751:4744]), .P(mul_out_593));
   mul8x8_wrap mul_594(.CLK(CLK), .W(W[4759:4752]), .IMG(IMG[4759:4752]), .P(mul_out_594));
   mul8x8_wrap mul_595(.CLK(CLK), .W(W[4767:4760]), .IMG(IMG[4767:4760]), .P(mul_out_595));
   mul8x8_wrap mul_596(.CLK(CLK), .W(W[4775:4768]), .IMG(IMG[4775:4768]), .P(mul_out_596));
   mul8x8_wrap mul_597(.CLK(CLK), .W(W[4783:4776]), .IMG(IMG[4783:4776]), .P(mul_out_597));
   mul8x8_wrap mul_598(.CLK(CLK), .W(W[4791:4784]), .IMG(IMG[4791:4784]), .P(mul_out_598));
   mul8x8_wrap mul_599(.CLK(CLK), .W(W[4799:4792]), .IMG(IMG[4799:4792]), .P(mul_out_599));
   mul8x8_wrap mul_600(.CLK(CLK), .W(W[4807:4800]), .IMG(IMG[4807:4800]), .P(mul_out_600));
   mul8x8_wrap mul_601(.CLK(CLK), .W(W[4815:4808]), .IMG(IMG[4815:4808]), .P(mul_out_601));
   mul8x8_wrap mul_602(.CLK(CLK), .W(W[4823:4816]), .IMG(IMG[4823:4816]), .P(mul_out_602));
   mul8x8_wrap mul_603(.CLK(CLK), .W(W[4831:4824]), .IMG(IMG[4831:4824]), .P(mul_out_603));
   mul8x8_wrap mul_604(.CLK(CLK), .W(W[4839:4832]), .IMG(IMG[4839:4832]), .P(mul_out_604));
   mul8x8_wrap mul_605(.CLK(CLK), .W(W[4847:4840]), .IMG(IMG[4847:4840]), .P(mul_out_605));
   mul8x8_wrap mul_606(.CLK(CLK), .W(W[4855:4848]), .IMG(IMG[4855:4848]), .P(mul_out_606));
   mul8x8_wrap mul_607(.CLK(CLK), .W(W[4863:4856]), .IMG(IMG[4863:4856]), .P(mul_out_607));
   mul8x8_wrap mul_608(.CLK(CLK), .W(W[4871:4864]), .IMG(IMG[4871:4864]), .P(mul_out_608));
   mul8x8_wrap mul_609(.CLK(CLK), .W(W[4879:4872]), .IMG(IMG[4879:4872]), .P(mul_out_609));
   mul8x8_wrap mul_610(.CLK(CLK), .W(W[4887:4880]), .IMG(IMG[4887:4880]), .P(mul_out_610));
   mul8x8_wrap mul_611(.CLK(CLK), .W(W[4895:4888]), .IMG(IMG[4895:4888]), .P(mul_out_611));
   mul8x8_wrap mul_612(.CLK(CLK), .W(W[4903:4896]), .IMG(IMG[4903:4896]), .P(mul_out_612));
   mul8x8_wrap mul_613(.CLK(CLK), .W(W[4911:4904]), .IMG(IMG[4911:4904]), .P(mul_out_613));
   mul8x8_wrap mul_614(.CLK(CLK), .W(W[4919:4912]), .IMG(IMG[4919:4912]), .P(mul_out_614));
   mul8x8_wrap mul_615(.CLK(CLK), .W(W[4927:4920]), .IMG(IMG[4927:4920]), .P(mul_out_615));
   mul8x8_wrap mul_616(.CLK(CLK), .W(W[4935:4928]), .IMG(IMG[4935:4928]), .P(mul_out_616));
   mul8x8_wrap mul_617(.CLK(CLK), .W(W[4943:4936]), .IMG(IMG[4943:4936]), .P(mul_out_617));
   mul8x8_wrap mul_618(.CLK(CLK), .W(W[4951:4944]), .IMG(IMG[4951:4944]), .P(mul_out_618));
   mul8x8_wrap mul_619(.CLK(CLK), .W(W[4959:4952]), .IMG(IMG[4959:4952]), .P(mul_out_619));
   mul8x8_wrap mul_620(.CLK(CLK), .W(W[4967:4960]), .IMG(IMG[4967:4960]), .P(mul_out_620));
   mul8x8_wrap mul_621(.CLK(CLK), .W(W[4975:4968]), .IMG(IMG[4975:4968]), .P(mul_out_621));
   mul8x8_wrap mul_622(.CLK(CLK), .W(W[4983:4976]), .IMG(IMG[4983:4976]), .P(mul_out_622));
   mul8x8_wrap mul_623(.CLK(CLK), .W(W[4991:4984]), .IMG(IMG[4991:4984]), .P(mul_out_623));
   mul8x8_wrap mul_624(.CLK(CLK), .W(W[4999:4992]), .IMG(IMG[4999:4992]), .P(mul_out_624));
   mul8x8_wrap mul_625(.CLK(CLK), .W(W[5007:5000]), .IMG(IMG[5007:5000]), .P(mul_out_625));
   mul8x8_wrap mul_626(.CLK(CLK), .W(W[5015:5008]), .IMG(IMG[5015:5008]), .P(mul_out_626));
   mul8x8_wrap mul_627(.CLK(CLK), .W(W[5023:5016]), .IMG(IMG[5023:5016]), .P(mul_out_627));
   mul8x8_wrap mul_628(.CLK(CLK), .W(W[5031:5024]), .IMG(IMG[5031:5024]), .P(mul_out_628));
   mul8x8_wrap mul_629(.CLK(CLK), .W(W[5039:5032]), .IMG(IMG[5039:5032]), .P(mul_out_629));
   mul8x8_wrap mul_630(.CLK(CLK), .W(W[5047:5040]), .IMG(IMG[5047:5040]), .P(mul_out_630));
   mul8x8_wrap mul_631(.CLK(CLK), .W(W[5055:5048]), .IMG(IMG[5055:5048]), .P(mul_out_631));
   mul8x8_wrap mul_632(.CLK(CLK), .W(W[5063:5056]), .IMG(IMG[5063:5056]), .P(mul_out_632));
   mul8x8_wrap mul_633(.CLK(CLK), .W(W[5071:5064]), .IMG(IMG[5071:5064]), .P(mul_out_633));
   mul8x8_wrap mul_634(.CLK(CLK), .W(W[5079:5072]), .IMG(IMG[5079:5072]), .P(mul_out_634));
   mul8x8_wrap mul_635(.CLK(CLK), .W(W[5087:5080]), .IMG(IMG[5087:5080]), .P(mul_out_635));
   mul8x8_wrap mul_636(.CLK(CLK), .W(W[5095:5088]), .IMG(IMG[5095:5088]), .P(mul_out_636));
   mul8x8_wrap mul_637(.CLK(CLK), .W(W[5103:5096]), .IMG(IMG[5103:5096]), .P(mul_out_637));
   mul8x8_wrap mul_638(.CLK(CLK), .W(W[5111:5104]), .IMG(IMG[5111:5104]), .P(mul_out_638));
   mul8x8_wrap mul_639(.CLK(CLK), .W(W[5119:5112]), .IMG(IMG[5119:5112]), .P(mul_out_639));
   mul8x8_wrap mul_640(.CLK(CLK), .W(W[5127:5120]), .IMG(IMG[5127:5120]), .P(mul_out_640));
   mul8x8_wrap mul_641(.CLK(CLK), .W(W[5135:5128]), .IMG(IMG[5135:5128]), .P(mul_out_641));
   mul8x8_wrap mul_642(.CLK(CLK), .W(W[5143:5136]), .IMG(IMG[5143:5136]), .P(mul_out_642));
   mul8x8_wrap mul_643(.CLK(CLK), .W(W[5151:5144]), .IMG(IMG[5151:5144]), .P(mul_out_643));
   mul8x8_wrap mul_644(.CLK(CLK), .W(W[5159:5152]), .IMG(IMG[5159:5152]), .P(mul_out_644));
   mul8x8_wrap mul_645(.CLK(CLK), .W(W[5167:5160]), .IMG(IMG[5167:5160]), .P(mul_out_645));
   mul8x8_wrap mul_646(.CLK(CLK), .W(W[5175:5168]), .IMG(IMG[5175:5168]), .P(mul_out_646));
   mul8x8_wrap mul_647(.CLK(CLK), .W(W[5183:5176]), .IMG(IMG[5183:5176]), .P(mul_out_647));
   mul8x8_wrap mul_648(.CLK(CLK), .W(W[5191:5184]), .IMG(IMG[5191:5184]), .P(mul_out_648));
   mul8x8_wrap mul_649(.CLK(CLK), .W(W[5199:5192]), .IMG(IMG[5199:5192]), .P(mul_out_649));
   mul8x8_wrap mul_650(.CLK(CLK), .W(W[5207:5200]), .IMG(IMG[5207:5200]), .P(mul_out_650));
   mul8x8_wrap mul_651(.CLK(CLK), .W(W[5215:5208]), .IMG(IMG[5215:5208]), .P(mul_out_651));
   mul8x8_wrap mul_652(.CLK(CLK), .W(W[5223:5216]), .IMG(IMG[5223:5216]), .P(mul_out_652));
   mul8x8_wrap mul_653(.CLK(CLK), .W(W[5231:5224]), .IMG(IMG[5231:5224]), .P(mul_out_653));
   mul8x8_wrap mul_654(.CLK(CLK), .W(W[5239:5232]), .IMG(IMG[5239:5232]), .P(mul_out_654));
   mul8x8_wrap mul_655(.CLK(CLK), .W(W[5247:5240]), .IMG(IMG[5247:5240]), .P(mul_out_655));
   mul8x8_wrap mul_656(.CLK(CLK), .W(W[5255:5248]), .IMG(IMG[5255:5248]), .P(mul_out_656));
   mul8x8_wrap mul_657(.CLK(CLK), .W(W[5263:5256]), .IMG(IMG[5263:5256]), .P(mul_out_657));
   mul8x8_wrap mul_658(.CLK(CLK), .W(W[5271:5264]), .IMG(IMG[5271:5264]), .P(mul_out_658));
   mul8x8_wrap mul_659(.CLK(CLK), .W(W[5279:5272]), .IMG(IMG[5279:5272]), .P(mul_out_659));
   mul8x8_wrap mul_660(.CLK(CLK), .W(W[5287:5280]), .IMG(IMG[5287:5280]), .P(mul_out_660));
   mul8x8_wrap mul_661(.CLK(CLK), .W(W[5295:5288]), .IMG(IMG[5295:5288]), .P(mul_out_661));
   mul8x8_wrap mul_662(.CLK(CLK), .W(W[5303:5296]), .IMG(IMG[5303:5296]), .P(mul_out_662));
   mul8x8_wrap mul_663(.CLK(CLK), .W(W[5311:5304]), .IMG(IMG[5311:5304]), .P(mul_out_663));
   mul8x8_wrap mul_664(.CLK(CLK), .W(W[5319:5312]), .IMG(IMG[5319:5312]), .P(mul_out_664));
   mul8x8_wrap mul_665(.CLK(CLK), .W(W[5327:5320]), .IMG(IMG[5327:5320]), .P(mul_out_665));
   mul8x8_wrap mul_666(.CLK(CLK), .W(W[5335:5328]), .IMG(IMG[5335:5328]), .P(mul_out_666));
   mul8x8_wrap mul_667(.CLK(CLK), .W(W[5343:5336]), .IMG(IMG[5343:5336]), .P(mul_out_667));
   mul8x8_wrap mul_668(.CLK(CLK), .W(W[5351:5344]), .IMG(IMG[5351:5344]), .P(mul_out_668));
   mul8x8_wrap mul_669(.CLK(CLK), .W(W[5359:5352]), .IMG(IMG[5359:5352]), .P(mul_out_669));
   mul8x8_wrap mul_670(.CLK(CLK), .W(W[5367:5360]), .IMG(IMG[5367:5360]), .P(mul_out_670));
   mul8x8_wrap mul_671(.CLK(CLK), .W(W[5375:5368]), .IMG(IMG[5375:5368]), .P(mul_out_671));
   mul8x8_wrap mul_672(.CLK(CLK), .W(W[5383:5376]), .IMG(IMG[5383:5376]), .P(mul_out_672));
   mul8x8_wrap mul_673(.CLK(CLK), .W(W[5391:5384]), .IMG(IMG[5391:5384]), .P(mul_out_673));
   mul8x8_wrap mul_674(.CLK(CLK), .W(W[5399:5392]), .IMG(IMG[5399:5392]), .P(mul_out_674));
   mul8x8_wrap mul_675(.CLK(CLK), .W(W[5407:5400]), .IMG(IMG[5407:5400]), .P(mul_out_675));
   mul8x8_wrap mul_676(.CLK(CLK), .W(W[5415:5408]), .IMG(IMG[5415:5408]), .P(mul_out_676));
   mul8x8_wrap mul_677(.CLK(CLK), .W(W[5423:5416]), .IMG(IMG[5423:5416]), .P(mul_out_677));
   mul8x8_wrap mul_678(.CLK(CLK), .W(W[5431:5424]), .IMG(IMG[5431:5424]), .P(mul_out_678));
   mul8x8_wrap mul_679(.CLK(CLK), .W(W[5439:5432]), .IMG(IMG[5439:5432]), .P(mul_out_679));
   mul8x8_wrap mul_680(.CLK(CLK), .W(W[5447:5440]), .IMG(IMG[5447:5440]), .P(mul_out_680));
   mul8x8_wrap mul_681(.CLK(CLK), .W(W[5455:5448]), .IMG(IMG[5455:5448]), .P(mul_out_681));
   mul8x8_wrap mul_682(.CLK(CLK), .W(W[5463:5456]), .IMG(IMG[5463:5456]), .P(mul_out_682));
   mul8x8_wrap mul_683(.CLK(CLK), .W(W[5471:5464]), .IMG(IMG[5471:5464]), .P(mul_out_683));
   mul8x8_wrap mul_684(.CLK(CLK), .W(W[5479:5472]), .IMG(IMG[5479:5472]), .P(mul_out_684));
   mul8x8_wrap mul_685(.CLK(CLK), .W(W[5487:5480]), .IMG(IMG[5487:5480]), .P(mul_out_685));
   mul8x8_wrap mul_686(.CLK(CLK), .W(W[5495:5488]), .IMG(IMG[5495:5488]), .P(mul_out_686));
   mul8x8_wrap mul_687(.CLK(CLK), .W(W[5503:5496]), .IMG(IMG[5503:5496]), .P(mul_out_687));
   mul8x8_wrap mul_688(.CLK(CLK), .W(W[5511:5504]), .IMG(IMG[5511:5504]), .P(mul_out_688));
   mul8x8_wrap mul_689(.CLK(CLK), .W(W[5519:5512]), .IMG(IMG[5519:5512]), .P(mul_out_689));
   mul8x8_wrap mul_690(.CLK(CLK), .W(W[5527:5520]), .IMG(IMG[5527:5520]), .P(mul_out_690));
   mul8x8_wrap mul_691(.CLK(CLK), .W(W[5535:5528]), .IMG(IMG[5535:5528]), .P(mul_out_691));
   mul8x8_wrap mul_692(.CLK(CLK), .W(W[5543:5536]), .IMG(IMG[5543:5536]), .P(mul_out_692));
   mul8x8_wrap mul_693(.CLK(CLK), .W(W[5551:5544]), .IMG(IMG[5551:5544]), .P(mul_out_693));
   mul8x8_wrap mul_694(.CLK(CLK), .W(W[5559:5552]), .IMG(IMG[5559:5552]), .P(mul_out_694));
   mul8x8_wrap mul_695(.CLK(CLK), .W(W[5567:5560]), .IMG(IMG[5567:5560]), .P(mul_out_695));
   mul8x8_wrap mul_696(.CLK(CLK), .W(W[5575:5568]), .IMG(IMG[5575:5568]), .P(mul_out_696));
   mul8x8_wrap mul_697(.CLK(CLK), .W(W[5583:5576]), .IMG(IMG[5583:5576]), .P(mul_out_697));
   mul8x8_wrap mul_698(.CLK(CLK), .W(W[5591:5584]), .IMG(IMG[5591:5584]), .P(mul_out_698));
   mul8x8_wrap mul_699(.CLK(CLK), .W(W[5599:5592]), .IMG(IMG[5599:5592]), .P(mul_out_699));
   mul8x8_wrap mul_700(.CLK(CLK), .W(W[5607:5600]), .IMG(IMG[5607:5600]), .P(mul_out_700));
   mul8x8_wrap mul_701(.CLK(CLK), .W(W[5615:5608]), .IMG(IMG[5615:5608]), .P(mul_out_701));
   mul8x8_wrap mul_702(.CLK(CLK), .W(W[5623:5616]), .IMG(IMG[5623:5616]), .P(mul_out_702));
   mul8x8_wrap mul_703(.CLK(CLK), .W(W[5631:5624]), .IMG(IMG[5631:5624]), .P(mul_out_703));
   mul8x8_wrap mul_704(.CLK(CLK), .W(W[5639:5632]), .IMG(IMG[5639:5632]), .P(mul_out_704));
   mul8x8_wrap mul_705(.CLK(CLK), .W(W[5647:5640]), .IMG(IMG[5647:5640]), .P(mul_out_705));
   mul8x8_wrap mul_706(.CLK(CLK), .W(W[5655:5648]), .IMG(IMG[5655:5648]), .P(mul_out_706));
   mul8x8_wrap mul_707(.CLK(CLK), .W(W[5663:5656]), .IMG(IMG[5663:5656]), .P(mul_out_707));
   mul8x8_wrap mul_708(.CLK(CLK), .W(W[5671:5664]), .IMG(IMG[5671:5664]), .P(mul_out_708));
   mul8x8_wrap mul_709(.CLK(CLK), .W(W[5679:5672]), .IMG(IMG[5679:5672]), .P(mul_out_709));
   mul8x8_wrap mul_710(.CLK(CLK), .W(W[5687:5680]), .IMG(IMG[5687:5680]), .P(mul_out_710));
   mul8x8_wrap mul_711(.CLK(CLK), .W(W[5695:5688]), .IMG(IMG[5695:5688]), .P(mul_out_711));
   mul8x8_wrap mul_712(.CLK(CLK), .W(W[5703:5696]), .IMG(IMG[5703:5696]), .P(mul_out_712));
   mul8x8_wrap mul_713(.CLK(CLK), .W(W[5711:5704]), .IMG(IMG[5711:5704]), .P(mul_out_713));
   mul8x8_wrap mul_714(.CLK(CLK), .W(W[5719:5712]), .IMG(IMG[5719:5712]), .P(mul_out_714));
   mul8x8_wrap mul_715(.CLK(CLK), .W(W[5727:5720]), .IMG(IMG[5727:5720]), .P(mul_out_715));
   mul8x8_wrap mul_716(.CLK(CLK), .W(W[5735:5728]), .IMG(IMG[5735:5728]), .P(mul_out_716));
   mul8x8_wrap mul_717(.CLK(CLK), .W(W[5743:5736]), .IMG(IMG[5743:5736]), .P(mul_out_717));
   mul8x8_wrap mul_718(.CLK(CLK), .W(W[5751:5744]), .IMG(IMG[5751:5744]), .P(mul_out_718));
   mul8x8_wrap mul_719(.CLK(CLK), .W(W[5759:5752]), .IMG(IMG[5759:5752]), .P(mul_out_719));
   mul8x8_wrap mul_720(.CLK(CLK), .W(W[5767:5760]), .IMG(IMG[5767:5760]), .P(mul_out_720));
   mul8x8_wrap mul_721(.CLK(CLK), .W(W[5775:5768]), .IMG(IMG[5775:5768]), .P(mul_out_721));
   mul8x8_wrap mul_722(.CLK(CLK), .W(W[5783:5776]), .IMG(IMG[5783:5776]), .P(mul_out_722));
   mul8x8_wrap mul_723(.CLK(CLK), .W(W[5791:5784]), .IMG(IMG[5791:5784]), .P(mul_out_723));
   mul8x8_wrap mul_724(.CLK(CLK), .W(W[5799:5792]), .IMG(IMG[5799:5792]), .P(mul_out_724));
   mul8x8_wrap mul_725(.CLK(CLK), .W(W[5807:5800]), .IMG(IMG[5807:5800]), .P(mul_out_725));
   mul8x8_wrap mul_726(.CLK(CLK), .W(W[5815:5808]), .IMG(IMG[5815:5808]), .P(mul_out_726));
   mul8x8_wrap mul_727(.CLK(CLK), .W(W[5823:5816]), .IMG(IMG[5823:5816]), .P(mul_out_727));
   mul8x8_wrap mul_728(.CLK(CLK), .W(W[5831:5824]), .IMG(IMG[5831:5824]), .P(mul_out_728));
   mul8x8_wrap mul_729(.CLK(CLK), .W(W[5839:5832]), .IMG(IMG[5839:5832]), .P(mul_out_729));
   mul8x8_wrap mul_730(.CLK(CLK), .W(W[5847:5840]), .IMG(IMG[5847:5840]), .P(mul_out_730));
   mul8x8_wrap mul_731(.CLK(CLK), .W(W[5855:5848]), .IMG(IMG[5855:5848]), .P(mul_out_731));
   mul8x8_wrap mul_732(.CLK(CLK), .W(W[5863:5856]), .IMG(IMG[5863:5856]), .P(mul_out_732));
   mul8x8_wrap mul_733(.CLK(CLK), .W(W[5871:5864]), .IMG(IMG[5871:5864]), .P(mul_out_733));
   mul8x8_wrap mul_734(.CLK(CLK), .W(W[5879:5872]), .IMG(IMG[5879:5872]), .P(mul_out_734));
   mul8x8_wrap mul_735(.CLK(CLK), .W(W[5887:5880]), .IMG(IMG[5887:5880]), .P(mul_out_735));
   mul8x8_wrap mul_736(.CLK(CLK), .W(W[5895:5888]), .IMG(IMG[5895:5888]), .P(mul_out_736));
   mul8x8_wrap mul_737(.CLK(CLK), .W(W[5903:5896]), .IMG(IMG[5903:5896]), .P(mul_out_737));
   mul8x8_wrap mul_738(.CLK(CLK), .W(W[5911:5904]), .IMG(IMG[5911:5904]), .P(mul_out_738));
   mul8x8_wrap mul_739(.CLK(CLK), .W(W[5919:5912]), .IMG(IMG[5919:5912]), .P(mul_out_739));
   mul8x8_wrap mul_740(.CLK(CLK), .W(W[5927:5920]), .IMG(IMG[5927:5920]), .P(mul_out_740));
   mul8x8_wrap mul_741(.CLK(CLK), .W(W[5935:5928]), .IMG(IMG[5935:5928]), .P(mul_out_741));
   mul8x8_wrap mul_742(.CLK(CLK), .W(W[5943:5936]), .IMG(IMG[5943:5936]), .P(mul_out_742));
   mul8x8_wrap mul_743(.CLK(CLK), .W(W[5951:5944]), .IMG(IMG[5951:5944]), .P(mul_out_743));
   mul8x8_wrap mul_744(.CLK(CLK), .W(W[5959:5952]), .IMG(IMG[5959:5952]), .P(mul_out_744));
   mul8x8_wrap mul_745(.CLK(CLK), .W(W[5967:5960]), .IMG(IMG[5967:5960]), .P(mul_out_745));
   mul8x8_wrap mul_746(.CLK(CLK), .W(W[5975:5968]), .IMG(IMG[5975:5968]), .P(mul_out_746));
   mul8x8_wrap mul_747(.CLK(CLK), .W(W[5983:5976]), .IMG(IMG[5983:5976]), .P(mul_out_747));
   mul8x8_wrap mul_748(.CLK(CLK), .W(W[5991:5984]), .IMG(IMG[5991:5984]), .P(mul_out_748));
   mul8x8_wrap mul_749(.CLK(CLK), .W(W[5999:5992]), .IMG(IMG[5999:5992]), .P(mul_out_749));
   mul8x8_wrap mul_750(.CLK(CLK), .W(W[6007:6000]), .IMG(IMG[6007:6000]), .P(mul_out_750));
   mul8x8_wrap mul_751(.CLK(CLK), .W(W[6015:6008]), .IMG(IMG[6015:6008]), .P(mul_out_751));
   mul8x8_wrap mul_752(.CLK(CLK), .W(W[6023:6016]), .IMG(IMG[6023:6016]), .P(mul_out_752));
   mul8x8_wrap mul_753(.CLK(CLK), .W(W[6031:6024]), .IMG(IMG[6031:6024]), .P(mul_out_753));
   mul8x8_wrap mul_754(.CLK(CLK), .W(W[6039:6032]), .IMG(IMG[6039:6032]), .P(mul_out_754));
   mul8x8_wrap mul_755(.CLK(CLK), .W(W[6047:6040]), .IMG(IMG[6047:6040]), .P(mul_out_755));
   mul8x8_wrap mul_756(.CLK(CLK), .W(W[6055:6048]), .IMG(IMG[6055:6048]), .P(mul_out_756));
   mul8x8_wrap mul_757(.CLK(CLK), .W(W[6063:6056]), .IMG(IMG[6063:6056]), .P(mul_out_757));
   mul8x8_wrap mul_758(.CLK(CLK), .W(W[6071:6064]), .IMG(IMG[6071:6064]), .P(mul_out_758));
   mul8x8_wrap mul_759(.CLK(CLK), .W(W[6079:6072]), .IMG(IMG[6079:6072]), .P(mul_out_759));
   mul8x8_wrap mul_760(.CLK(CLK), .W(W[6087:6080]), .IMG(IMG[6087:6080]), .P(mul_out_760));
   mul8x8_wrap mul_761(.CLK(CLK), .W(W[6095:6088]), .IMG(IMG[6095:6088]), .P(mul_out_761));
   mul8x8_wrap mul_762(.CLK(CLK), .W(W[6103:6096]), .IMG(IMG[6103:6096]), .P(mul_out_762));
   mul8x8_wrap mul_763(.CLK(CLK), .W(W[6111:6104]), .IMG(IMG[6111:6104]), .P(mul_out_763));
   mul8x8_wrap mul_764(.CLK(CLK), .W(W[6119:6112]), .IMG(IMG[6119:6112]), .P(mul_out_764));
   mul8x8_wrap mul_765(.CLK(CLK), .W(W[6127:6120]), .IMG(IMG[6127:6120]), .P(mul_out_765));
   mul8x8_wrap mul_766(.CLK(CLK), .W(W[6135:6128]), .IMG(IMG[6135:6128]), .P(mul_out_766));
   mul8x8_wrap mul_767(.CLK(CLK), .W(W[6143:6136]), .IMG(IMG[6143:6136]), .P(mul_out_767));
   mul8x8_wrap mul_768(.CLK(CLK), .W(W[6151:6144]), .IMG(IMG[6151:6144]), .P(mul_out_768));
   mul8x8_wrap mul_769(.CLK(CLK), .W(W[6159:6152]), .IMG(IMG[6159:6152]), .P(mul_out_769));
   mul8x8_wrap mul_770(.CLK(CLK), .W(W[6167:6160]), .IMG(IMG[6167:6160]), .P(mul_out_770));
   mul8x8_wrap mul_771(.CLK(CLK), .W(W[6175:6168]), .IMG(IMG[6175:6168]), .P(mul_out_771));
   mul8x8_wrap mul_772(.CLK(CLK), .W(W[6183:6176]), .IMG(IMG[6183:6176]), .P(mul_out_772));
   mul8x8_wrap mul_773(.CLK(CLK), .W(W[6191:6184]), .IMG(IMG[6191:6184]), .P(mul_out_773));
   mul8x8_wrap mul_774(.CLK(CLK), .W(W[6199:6192]), .IMG(IMG[6199:6192]), .P(mul_out_774));
   mul8x8_wrap mul_775(.CLK(CLK), .W(W[6207:6200]), .IMG(IMG[6207:6200]), .P(mul_out_775));
   mul8x8_wrap mul_776(.CLK(CLK), .W(W[6215:6208]), .IMG(IMG[6215:6208]), .P(mul_out_776));
   mul8x8_wrap mul_777(.CLK(CLK), .W(W[6223:6216]), .IMG(IMG[6223:6216]), .P(mul_out_777));
   mul8x8_wrap mul_778(.CLK(CLK), .W(W[6231:6224]), .IMG(IMG[6231:6224]), .P(mul_out_778));
   mul8x8_wrap mul_779(.CLK(CLK), .W(W[6239:6232]), .IMG(IMG[6239:6232]), .P(mul_out_779));
   mul8x8_wrap mul_780(.CLK(CLK), .W(W[6247:6240]), .IMG(IMG[6247:6240]), .P(mul_out_780));
   mul8x8_wrap mul_781(.CLK(CLK), .W(W[6255:6248]), .IMG(IMG[6255:6248]), .P(mul_out_781));
   mul8x8_wrap mul_782(.CLK(CLK), .W(W[6263:6256]), .IMG(IMG[6263:6256]), .P(mul_out_782));
   mul8x8_wrap mul_783(.CLK(CLK), .W(W[6271:6264]), .IMG(IMG[6271:6264]), .P(mul_out_783));

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_00 <= 0;
      end else begin
	 add_00 <= mul_out_0 + mul_out_1 + mul_out_2 + mul_out_3 + mul_out_4 + mul_out_5 + mul_out_6 + mul_out_7 + mul_out_8 + mul_out_9 + mul_out_10 + mul_out_11 + mul_out_12 + mul_out_13 + mul_out_14 + mul_out_15 + mul_out_16 + mul_out_17 + mul_out_18 + mul_out_19 + mul_out_20 + mul_out_21 + mul_out_22 + mul_out_23 + mul_out_24 + mul_out_25 + mul_out_26 + mul_out_27;
      end
   end


   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_01 <= 0;
      end else begin
	 add_01 <= mul_out_28 + mul_out_29 + mul_out_30 + mul_out_31 + mul_out_32 + mul_out_33 + mul_out_34 + mul_out_35 + mul_out_36 + mul_out_37 + mul_out_38 + mul_out_39 + mul_out_40 + mul_out_41 + mul_out_42 + mul_out_43 + mul_out_44 + mul_out_45 + mul_out_46 + mul_out_47 + mul_out_48 + mul_out_49 + mul_out_50 + mul_out_51 + mul_out_52 + mul_out_53 + mul_out_54 + mul_out_55;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_02 <= 0;
      end else begin
	 add_02 <= mul_out_56 + mul_out_57 + mul_out_58 + mul_out_59 + mul_out_60 + mul_out_61 + mul_out_62 + mul_out_63 + mul_out_64 + mul_out_65 + mul_out_66 + mul_out_67 + mul_out_68 + mul_out_69 + mul_out_70 + mul_out_71 + mul_out_72 + mul_out_73 + mul_out_74 + mul_out_75 + mul_out_76 + mul_out_77 + mul_out_78 + mul_out_79 + mul_out_80 + mul_out_81 + mul_out_82 + mul_out_83;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_03 <= 0;
      end else begin
	 add_03 <= mul_out_84 + mul_out_85 + mul_out_86 + mul_out_87 + mul_out_88 + mul_out_89 + mul_out_90 + mul_out_91 + mul_out_92 + mul_out_93 + mul_out_94 + mul_out_95 + mul_out_96 + mul_out_97 + mul_out_98 + mul_out_99 + mul_out_100 + mul_out_101 + mul_out_102 + mul_out_103 + mul_out_104 + mul_out_105 + mul_out_106 + mul_out_107 + mul_out_108 + mul_out_109 + mul_out_110 + mul_out_111;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_04 <= 0;
      end else begin
	 add_04 <= mul_out_112 + mul_out_113 + mul_out_114 + mul_out_115 + mul_out_116 + mul_out_117 + mul_out_118 + mul_out_119 + mul_out_120 + mul_out_121 + mul_out_122 + mul_out_123 + mul_out_124 + mul_out_125 + mul_out_126 + mul_out_127 + mul_out_128 + mul_out_129 + mul_out_130 + mul_out_131 + mul_out_132 + mul_out_133 + mul_out_134 + mul_out_135 + mul_out_136 + mul_out_137 + mul_out_138 + mul_out_139;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_05 <= 0;
      end else begin
	 add_05 <= mul_out_140 + mul_out_141 + mul_out_142 + mul_out_143 + mul_out_144 + mul_out_145 + mul_out_146 + mul_out_147 + mul_out_148 + mul_out_149 + mul_out_150 + mul_out_151 + mul_out_152 + mul_out_153 + mul_out_154 + mul_out_155 + mul_out_156 + mul_out_157 + mul_out_158 + mul_out_159 + mul_out_160 + mul_out_161 + mul_out_162 + mul_out_163 + mul_out_164 + mul_out_165 + mul_out_166 + mul_out_167;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_06 <= 0;
      end else begin
	 add_06 <= mul_out_168 + mul_out_169 + mul_out_170 + mul_out_171 + mul_out_172 + mul_out_173 + mul_out_174 + mul_out_175 + mul_out_176 + mul_out_177 + mul_out_178 + mul_out_179 + mul_out_180 + mul_out_181 + mul_out_182 + mul_out_183 + mul_out_184 + mul_out_185 + mul_out_186 + mul_out_187 + mul_out_188 + mul_out_189 + mul_out_190 + mul_out_191 + mul_out_192 + mul_out_193 + mul_out_194 + mul_out_195;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_07 <= 0;
      end else begin
	 add_07 <= mul_out_196 + mul_out_197 + mul_out_198 + mul_out_199 + mul_out_200 + mul_out_201 + mul_out_202 + mul_out_203 + mul_out_204 + mul_out_205 + mul_out_206 + mul_out_207 + mul_out_208 + mul_out_209 + mul_out_210 + mul_out_211 + mul_out_212 + mul_out_213 + mul_out_214 + mul_out_215 + mul_out_216 + mul_out_217 + mul_out_218 + mul_out_219 + mul_out_220 + mul_out_221 + mul_out_222 + mul_out_223;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_08 <= 0;
      end else begin
	 add_08 <= mul_out_224 + mul_out_225 + mul_out_226 + mul_out_227 + mul_out_228 + mul_out_229 + mul_out_230 + mul_out_231 + mul_out_232 + mul_out_233 + mul_out_234 + mul_out_235 + mul_out_236 + mul_out_237 + mul_out_238 + mul_out_239 + mul_out_240 + mul_out_241 + mul_out_242 + mul_out_243 + mul_out_244 + mul_out_245 + mul_out_246 + mul_out_247 + mul_out_248 + mul_out_249 + mul_out_250 + mul_out_251;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_09 <= 0;
      end else begin
	 add_09 <= mul_out_252 + mul_out_253 + mul_out_254 + mul_out_255 + mul_out_256 + mul_out_257 + mul_out_258 + mul_out_259 + mul_out_260 + mul_out_261 + mul_out_262 + mul_out_263 + mul_out_264 + mul_out_265 + mul_out_266 + mul_out_267 + mul_out_268 + mul_out_269 + mul_out_270 + mul_out_271 + mul_out_272 + mul_out_273 + mul_out_274 + mul_out_275 + mul_out_276 + mul_out_277 + mul_out_278 + mul_out_279;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_10 <= 0;
      end else begin
	 add_10 <= mul_out_280 + mul_out_281 + mul_out_282 + mul_out_283 + mul_out_284 + mul_out_285 + mul_out_286 + mul_out_287 + mul_out_288 + mul_out_289 + mul_out_290 + mul_out_291 + mul_out_292 + mul_out_293 + mul_out_294 + mul_out_295 + mul_out_296 + mul_out_297 + mul_out_298 + mul_out_299 + mul_out_300 + mul_out_301 + mul_out_302 + mul_out_303 + mul_out_304 + mul_out_305 + mul_out_306 + mul_out_307;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_11 <= 0;
      end else begin
	 add_11 <= mul_out_308 + mul_out_309 + mul_out_310 + mul_out_311 + mul_out_312 + mul_out_313 + mul_out_314 + mul_out_315 + mul_out_316 + mul_out_317 + mul_out_318 + mul_out_319 + mul_out_320 + mul_out_321 + mul_out_322 + mul_out_323 + mul_out_324 + mul_out_325 + mul_out_326 + mul_out_327 + mul_out_328 + mul_out_329 + mul_out_330 + mul_out_331 + mul_out_332 + mul_out_333 + mul_out_334 + mul_out_335;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_12 <= 0;
      end else begin
	 add_12 <= mul_out_336 + mul_out_337 + mul_out_338 + mul_out_339 + mul_out_340 + mul_out_341 + mul_out_342 + mul_out_343 + mul_out_344 + mul_out_345 + mul_out_346 + mul_out_347 + mul_out_348 + mul_out_349 + mul_out_350 + mul_out_351 + mul_out_352 + mul_out_353 + mul_out_354 + mul_out_355 + mul_out_356 + mul_out_357 + mul_out_358 + mul_out_359 + mul_out_360 + mul_out_361 + mul_out_362 + mul_out_363;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_13 <= 0;
      end else begin
	 add_13 <= mul_out_364 + mul_out_365 + mul_out_366 + mul_out_367 + mul_out_368 + mul_out_369 + mul_out_370 + mul_out_371 + mul_out_372 + mul_out_373 + mul_out_374 + mul_out_375 + mul_out_376 + mul_out_377 + mul_out_378 + mul_out_379 + mul_out_380 + mul_out_381 + mul_out_382 + mul_out_383 + mul_out_384 + mul_out_385 + mul_out_386 + mul_out_387 + mul_out_388 + mul_out_389 + mul_out_390 + mul_out_391;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_14 <= 0;
      end else begin
	 add_14 <= mul_out_392 + mul_out_393 + mul_out_394 + mul_out_395 + mul_out_396 + mul_out_397 + mul_out_398 + mul_out_399 + mul_out_400 + mul_out_401 + mul_out_402 + mul_out_403 + mul_out_404 + mul_out_405 + mul_out_406 + mul_out_407 + mul_out_408 + mul_out_409 + mul_out_410 + mul_out_411 + mul_out_412 + mul_out_413 + mul_out_414 + mul_out_415 + mul_out_416 + mul_out_417 + mul_out_418 + mul_out_419;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_15 <= 0;
      end else begin
	 add_15 <= mul_out_420 + mul_out_421 + mul_out_422 + mul_out_423 + mul_out_424 + mul_out_425 + mul_out_426 + mul_out_427 + mul_out_428 + mul_out_429 + mul_out_430 + mul_out_431 + mul_out_432 + mul_out_433 + mul_out_434 + mul_out_435 + mul_out_436 + mul_out_437 + mul_out_438 + mul_out_439 + mul_out_440 + mul_out_441 + mul_out_442 + mul_out_443 + mul_out_444 + mul_out_445 + mul_out_446 + mul_out_447;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_16 <= 0;
      end else begin
	 add_16 <= mul_out_448 + mul_out_449 + mul_out_450 + mul_out_451 + mul_out_452 + mul_out_453 + mul_out_454 + mul_out_455 + mul_out_456 + mul_out_457 + mul_out_458 + mul_out_459 + mul_out_460 + mul_out_461 + mul_out_462 + mul_out_463 + mul_out_464 + mul_out_465 + mul_out_466 + mul_out_467 + mul_out_468 + mul_out_469 + mul_out_470 + mul_out_471 + mul_out_472 + mul_out_473 + mul_out_474 + mul_out_475;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_17 <= 0;
      end else begin
	 add_17 <= mul_out_476 + mul_out_477 + mul_out_478 + mul_out_479 + mul_out_480 + mul_out_481 + mul_out_482 + mul_out_483 + mul_out_484 + mul_out_485 + mul_out_486 + mul_out_487 + mul_out_488 + mul_out_489 + mul_out_490 + mul_out_491 + mul_out_492 + mul_out_493 + mul_out_494 + mul_out_495 + mul_out_496 + mul_out_497 + mul_out_498 + mul_out_499 + mul_out_500 + mul_out_501 + mul_out_502 + mul_out_503;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_18 <= 0;
      end else begin
	 add_18 <= mul_out_504 + mul_out_505 + mul_out_506 + mul_out_507 + mul_out_508 + mul_out_509 + mul_out_510 + mul_out_511 + mul_out_512 + mul_out_513 + mul_out_514 + mul_out_515 + mul_out_516 + mul_out_517 + mul_out_518 + mul_out_519 + mul_out_520 + mul_out_521 + mul_out_522 + mul_out_523 + mul_out_524 + mul_out_525 + mul_out_526 + mul_out_527 + mul_out_528 + mul_out_529 + mul_out_530 + mul_out_531;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_19 <= 0;
      end else begin
	 add_19 <= mul_out_532 + mul_out_533 + mul_out_534 + mul_out_535 + mul_out_536 + mul_out_537 + mul_out_538 + mul_out_539 + mul_out_540 + mul_out_541 + mul_out_542 + mul_out_543 + mul_out_544 + mul_out_545 + mul_out_546 + mul_out_547 + mul_out_548 + mul_out_549 + mul_out_550 + mul_out_551 + mul_out_552 + mul_out_553 + mul_out_554 + mul_out_555 + mul_out_556 + mul_out_557 + mul_out_558 + mul_out_559;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_20 <= 0;
      end else begin
	 add_20 <= mul_out_560 + mul_out_561 + mul_out_562 + mul_out_563 + mul_out_564 + mul_out_565 + mul_out_566 + mul_out_567 + mul_out_568 + mul_out_569 + mul_out_570 + mul_out_571 + mul_out_572 + mul_out_573 + mul_out_574 + mul_out_575 + mul_out_576 + mul_out_577 + mul_out_578 + mul_out_579 + mul_out_580 + mul_out_581 + mul_out_582 + mul_out_583 + mul_out_584 + mul_out_585 + mul_out_586 + mul_out_587;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_21 <= 0;
      end else begin
	 add_21 <= mul_out_588 + mul_out_589 + mul_out_590 + mul_out_591 + mul_out_592 + mul_out_593 + mul_out_594 + mul_out_595 + mul_out_596 + mul_out_597 + mul_out_598 + mul_out_599 + mul_out_600 + mul_out_601 + mul_out_602 + mul_out_603 + mul_out_604 + mul_out_605 + mul_out_606 + mul_out_607 + mul_out_608 + mul_out_609 + mul_out_610 + mul_out_611 + mul_out_612 + mul_out_613 + mul_out_614 + mul_out_615;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_22 <= 0;
      end else begin
	 add_22 <= mul_out_616 + mul_out_617 + mul_out_618 + mul_out_619 + mul_out_620 + mul_out_621 + mul_out_622 + mul_out_623 + mul_out_624 + mul_out_625 + mul_out_626 + mul_out_627 + mul_out_628 + mul_out_629 + mul_out_630 + mul_out_631 + mul_out_632 + mul_out_633 + mul_out_634 + mul_out_635 + mul_out_636 + mul_out_637 + mul_out_638 + mul_out_639 + mul_out_640 + mul_out_641 + mul_out_642 + mul_out_643;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_23 <= 0;
      end else begin
	 add_23 <= mul_out_644 + mul_out_645 + mul_out_646 + mul_out_647 + mul_out_648 + mul_out_649 + mul_out_650 + mul_out_651 + mul_out_652 + mul_out_653 + mul_out_654 + mul_out_655 + mul_out_656 + mul_out_657 + mul_out_658 + mul_out_659 + mul_out_660 + mul_out_661 + mul_out_662 + mul_out_663 + mul_out_664 + mul_out_665 + mul_out_666 + mul_out_667 + mul_out_668 + mul_out_669 + mul_out_670 + mul_out_671;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_24 <= 0;
      end else begin
	 add_24 <= mul_out_672 + mul_out_673 + mul_out_674 + mul_out_675 + mul_out_676 + mul_out_677 + mul_out_678 + mul_out_679 + mul_out_680 + mul_out_681 + mul_out_682 + mul_out_683 + mul_out_684 + mul_out_685 + mul_out_686 + mul_out_687 + mul_out_688 + mul_out_689 + mul_out_690 + mul_out_691 + mul_out_692 + mul_out_693 + mul_out_694 + mul_out_695 + mul_out_696 + mul_out_697 + mul_out_698 + mul_out_699;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_25 <= 0;
      end else begin
	 add_25 <= mul_out_700 + mul_out_701 + mul_out_702 + mul_out_703 + mul_out_704 + mul_out_705 + mul_out_706 + mul_out_707 + mul_out_708 + mul_out_709 + mul_out_710 + mul_out_711 + mul_out_712 + mul_out_713 + mul_out_714 + mul_out_715 + mul_out_716 + mul_out_717 + mul_out_718 + mul_out_719 + mul_out_720 + mul_out_721 + mul_out_722 + mul_out_723 + mul_out_724 + mul_out_725 + mul_out_726 + mul_out_727;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_26 <= 0;
      end else begin
	 add_26 <= mul_out_728 + mul_out_729 + mul_out_730 + mul_out_731 + mul_out_732 + mul_out_733 + mul_out_734 + mul_out_735 + mul_out_736 + mul_out_737 + mul_out_738 + mul_out_739 + mul_out_740 + mul_out_741 + mul_out_742 + mul_out_743 + mul_out_744 + mul_out_745 + mul_out_746 + mul_out_747 + mul_out_748 + mul_out_749 + mul_out_750 + mul_out_751 + mul_out_752 + mul_out_753 + mul_out_754 + mul_out_755;
      end
   end

   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 add_27 <= 0;
      end else begin
	 add_27 <= mul_out_756 + mul_out_757 + mul_out_758 + mul_out_759 + mul_out_760 + mul_out_761 + mul_out_762 + mul_out_763 + mul_out_764 + mul_out_765 + mul_out_766 + mul_out_767 + mul_out_768 + mul_out_769 + mul_out_770 + mul_out_771 + mul_out_772 + mul_out_773 + mul_out_774 + mul_out_775 + mul_out_776 + mul_out_777 + mul_out_778 + mul_out_779 + mul_out_780 + mul_out_781 + mul_out_782 + mul_out_783;
      end
   end


   always @ (posedge CLK or negedge RESET_X)begin
      if(RESET_X == 0)begin
	 RESULT <= 0;
      end else begin
	 RESULT <= add_00 + add_01 + add_02 + add_03 + add_04 + add_05 + add_06 + add_07 + add_08 + add_09 +
		   add_10 + add_11 + add_12 + add_13 + add_14 + add_15 + add_16 + add_17 + add_18 + add_19 +
		   add_20 + add_21 + add_22 + add_23 + add_24 + add_25 + add_26 + add_27 + B;
	 
      end
   end



endmodule // mul_add_core
