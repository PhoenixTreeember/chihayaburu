module softmax_top
  (
   input 	 CLK,
   input 	 RESET_X,
   input 	 WR,
   input 	 RD,
   input [17:0]  ADR,
   input [31:0]  WDATA,
   output [31:0] RDATA   
   );


   

endmodule // softmax_top
